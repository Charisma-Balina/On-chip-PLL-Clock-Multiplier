* SKY130 Spice File.
.param  globalk=1
.param  localkswitch=1
.param  capunits = '1.0*1e-6'
.param
+ mcp1f_ca_w_0_150_s_0_210 = 8.04e-05  mcp1f_cc_w_0_150_s_0_210 = 6.56e-11  mcp1f_cf_w_0_150_s_0_210 = 8.68e-12
+ mcp1f_ca_w_0_150_s_0_263 = 8.04e-05  mcp1f_cc_w_0_150_s_0_263 = 5.50e-11  mcp1f_cf_w_0_150_s_0_263 = 1.04e-11
+ mcp1f_ca_w_0_150_s_0_315 = 8.04e-05  mcp1f_cc_w_0_150_s_0_315 = 4.79e-11  mcp1f_cf_w_0_150_s_0_315 = 1.20e-11
+ mcp1f_ca_w_0_150_s_0_420 = 8.04e-05  mcp1f_cc_w_0_150_s_0_420 = 3.77e-11  mcp1f_cf_w_0_150_s_0_420 = 1.52e-11
+ mcp1f_ca_w_0_150_s_0_525 = 8.04e-05  mcp1f_cc_w_0_150_s_0_525 = 3.13e-11  mcp1f_cf_w_0_150_s_0_525 = 1.79e-11
+ mcp1f_ca_w_0_150_s_0_630 = 8.04e-05  mcp1f_cc_w_0_150_s_0_630 = 2.67e-11  mcp1f_cf_w_0_150_s_0_630 = 2.03e-11
+ mcp1f_ca_w_0_150_s_0_840 = 8.04e-05  mcp1f_cc_w_0_150_s_0_840 = 2.01e-11  mcp1f_cf_w_0_150_s_0_840 = 2.45e-11
+ mcp1f_ca_w_0_150_s_1_260 = 8.04e-05  mcp1f_cc_w_0_150_s_1_260 = 1.21e-11  mcp1f_cf_w_0_150_s_1_260 = 3.07e-11
+ mcp1f_ca_w_0_150_s_2_310 = 8.04e-05  mcp1f_cc_w_0_150_s_2_310 = 5.38e-12  mcp1f_cf_w_0_150_s_2_310 = 3.68e-11
+ mcp1f_ca_w_0_150_s_5_250 = 8.04e-05  mcp1f_cc_w_0_150_s_5_250 = 1.25e-12  mcp1f_cf_w_0_150_s_5_250 = 4.09e-11
+ mcp1f_ca_w_1_200_s_0_210 = 8.04e-05  mcp1f_cc_w_1_200_s_0_210 = 8.41e-11  mcp1f_cf_w_1_200_s_0_210 = 8.62e-12
+ mcp1f_ca_w_1_200_s_0_263 = 8.04e-05  mcp1f_cc_w_1_200_s_0_263 = 7.22e-11  mcp1f_cf_w_1_200_s_0_263 = 1.04e-11
+ mcp1f_ca_w_1_200_s_0_315 = 8.04e-05  mcp1f_cc_w_1_200_s_0_315 = 6.38e-11  mcp1f_cf_w_1_200_s_0_315 = 1.20e-11
+ mcp1f_ca_w_1_200_s_0_420 = 8.04e-05  mcp1f_cc_w_1_200_s_0_420 = 5.24e-11  mcp1f_cf_w_1_200_s_0_420 = 1.52e-11
+ mcp1f_ca_w_1_200_s_0_525 = 8.04e-05  mcp1f_cc_w_1_200_s_0_525 = 4.46e-11  mcp1f_cf_w_1_200_s_0_525 = 1.80e-11
+ mcp1f_ca_w_1_200_s_0_630 = 8.04e-05  mcp1f_cc_w_1_200_s_0_630 = 3.89e-11  mcp1f_cf_w_1_200_s_0_630 = 2.06e-11
+ mcp1f_ca_w_1_200_s_0_840 = 8.04e-05  mcp1f_cc_w_1_200_s_0_840 = 3.10e-11  mcp1f_cf_w_1_200_s_0_840 = 2.51e-11
+ mcp1f_ca_w_1_200_s_1_260 = 8.04e-05  mcp1f_cc_w_1_200_s_1_260 = 2.16e-11  mcp1f_cf_w_1_200_s_1_260 = 3.17e-11
+ mcp1f_ca_w_1_200_s_2_310 = 8.04e-05  mcp1f_cc_w_1_200_s_2_310 = 1.11e-11  mcp1f_cf_w_1_200_s_2_310 = 4.07e-11
+ mcp1f_ca_w_1_200_s_5_250 = 8.04e-05  mcp1f_cc_w_1_200_s_5_250 = 3.60e-12  mcp1f_cf_w_1_200_s_5_250 = 4.80e-11
+ mcl1f_ca_w_0_170_s_0_180 = 2.93e-05  mcl1f_cc_w_0_170_s_0_180 = 6.50e-11  mcl1f_cf_w_0_170_s_0_180 = 3.07e-12
+ mcl1f_ca_w_0_170_s_0_225 = 2.93e-05  mcl1f_cc_w_0_170_s_0_225 = 5.73e-11  mcl1f_cf_w_0_170_s_0_225 = 3.70e-12
+ mcl1f_ca_w_0_170_s_0_270 = 2.93e-05  mcl1f_cc_w_0_170_s_0_270 = 5.22e-11  mcl1f_cf_w_0_170_s_0_270 = 4.31e-12
+ mcl1f_ca_w_0_170_s_0_360 = 2.93e-05  mcl1f_cc_w_0_170_s_0_360 = 4.39e-11  mcl1f_cf_w_0_170_s_0_360 = 5.67e-12
+ mcl1f_ca_w_0_170_s_0_450 = 2.93e-05  mcl1f_cc_w_0_170_s_0_450 = 3.89e-11  mcl1f_cf_w_0_170_s_0_450 = 6.66e-12
+ mcl1f_ca_w_0_170_s_0_540 = 2.93e-05  mcl1f_cc_w_0_170_s_0_540 = 3.44e-11  mcl1f_cf_w_0_170_s_0_540 = 8.00e-12
+ mcl1f_ca_w_0_170_s_0_720 = 2.93e-05  mcl1f_cc_w_0_170_s_0_720 = 2.84e-11  mcl1f_cf_w_0_170_s_0_720 = 1.01e-11
+ mcl1f_ca_w_0_170_s_1_080 = 2.93e-05  mcl1f_cc_w_0_170_s_1_080 = 2.09e-11  mcl1f_cf_w_0_170_s_1_080 = 1.39e-11
+ mcl1f_ca_w_0_170_s_1_980 = 2.93e-05  mcl1f_cc_w_0_170_s_1_980 = 1.19e-11  mcl1f_cf_w_0_170_s_1_980 = 2.00e-11
+ mcl1f_ca_w_0_170_s_4_500 = 2.93e-05  mcl1f_cc_w_0_170_s_4_500 = 3.88e-12  mcl1f_cf_w_0_170_s_4_500 = 2.71e-11
+ mcl1f_ca_w_1_360_s_0_180 = 2.93e-05  mcl1f_cc_w_1_360_s_0_180 = 8.88e-11  mcl1f_cf_w_1_360_s_0_180 = 3.07e-12
+ mcl1f_ca_w_1_360_s_0_225 = 2.93e-05  mcl1f_cc_w_1_360_s_0_225 = 7.97e-11  mcl1f_cf_w_1_360_s_0_225 = 3.70e-12
+ mcl1f_ca_w_1_360_s_0_270 = 2.93e-05  mcl1f_cc_w_1_360_s_0_270 = 7.29e-11  mcl1f_cf_w_1_360_s_0_270 = 4.32e-12
+ mcl1f_ca_w_1_360_s_0_360 = 2.93e-05  mcl1f_cc_w_1_360_s_0_360 = 6.29e-11  mcl1f_cf_w_1_360_s_0_360 = 5.54e-12
+ mcl1f_ca_w_1_360_s_0_450 = 2.93e-05  mcl1f_cc_w_1_360_s_0_450 = 5.59e-11  mcl1f_cf_w_1_360_s_0_450 = 6.73e-12
+ mcl1f_ca_w_1_360_s_0_540 = 2.93e-05  mcl1f_cc_w_1_360_s_0_540 = 5.05e-11  mcl1f_cf_w_1_360_s_0_540 = 7.88e-12
+ mcl1f_ca_w_1_360_s_0_720 = 2.93e-05  mcl1f_cc_w_1_360_s_0_720 = 4.26e-11  mcl1f_cf_w_1_360_s_0_720 = 1.01e-11
+ mcl1f_ca_w_1_360_s_1_080 = 2.93e-05  mcl1f_cc_w_1_360_s_1_080 = 3.28e-11  mcl1f_cf_w_1_360_s_1_080 = 1.40e-11
+ mcl1f_ca_w_1_360_s_1_980 = 2.93e-05  mcl1f_cc_w_1_360_s_1_980 = 2.02e-11  mcl1f_cf_w_1_360_s_1_980 = 2.17e-11
+ mcl1f_ca_w_1_360_s_4_500 = 2.93e-05  mcl1f_cc_w_1_360_s_4_500 = 7.90e-12  mcl1f_cf_w_1_360_s_4_500 = 3.19e-11
+ mcl1d_ca_w_0_170_s_0_180 = 4.53e-05  mcl1d_cc_w_0_170_s_0_180 = 6.28e-11  mcl1d_cf_w_0_170_s_0_180 = 4.69e-12
+ mcl1d_ca_w_0_170_s_0_225 = 4.53e-05  mcl1d_cc_w_0_170_s_0_225 = 5.50e-11  mcl1d_cf_w_0_170_s_0_225 = 5.62e-12
+ mcl1d_ca_w_0_170_s_0_270 = 4.53e-05  mcl1d_cc_w_0_170_s_0_270 = 4.97e-11  mcl1d_cf_w_0_170_s_0_270 = 6.52e-12
+ mcl1d_ca_w_0_170_s_0_360 = 4.53e-05  mcl1d_cc_w_0_170_s_0_360 = 4.11e-11  mcl1d_cf_w_0_170_s_0_360 = 8.52e-12
+ mcl1d_ca_w_0_170_s_0_450 = 4.53e-05  mcl1d_cc_w_0_170_s_0_450 = 3.58e-11  mcl1d_cf_w_0_170_s_0_450 = 9.96e-12
+ mcl1d_ca_w_0_170_s_0_540 = 4.53e-05  mcl1d_cc_w_0_170_s_0_540 = 3.11e-11  mcl1d_cf_w_0_170_s_0_540 = 1.18e-11
+ mcl1d_ca_w_0_170_s_0_720 = 4.53e-05  mcl1d_cc_w_0_170_s_0_720 = 2.48e-11  mcl1d_cf_w_0_170_s_0_720 = 1.48e-11
+ mcl1d_ca_w_0_170_s_1_080 = 4.53e-05  mcl1d_cc_w_0_170_s_1_080 = 1.71e-11  mcl1d_cf_w_0_170_s_1_080 = 1.95e-11
+ mcl1d_ca_w_0_170_s_1_980 = 4.53e-05  mcl1d_cc_w_0_170_s_1_980 = 8.68e-12  mcl1d_cf_w_0_170_s_1_980 = 2.62e-11
+ mcl1d_ca_w_0_170_s_4_500 = 4.53e-05  mcl1d_cc_w_0_170_s_4_500 = 2.47e-12  mcl1d_cf_w_0_170_s_4_500 = 3.21e-11
+ mcl1d_ca_w_1_360_s_0_180 = 4.53e-05  mcl1d_cc_w_1_360_s_0_180 = 8.41e-11  mcl1d_cf_w_1_360_s_0_180 = 4.69e-12
+ mcl1d_ca_w_1_360_s_0_225 = 4.53e-05  mcl1d_cc_w_1_360_s_0_225 = 7.51e-11  mcl1d_cf_w_1_360_s_0_225 = 5.63e-12
+ mcl1d_ca_w_1_360_s_0_270 = 4.53e-05  mcl1d_cc_w_1_360_s_0_270 = 6.82e-11  mcl1d_cf_w_1_360_s_0_270 = 6.56e-12
+ mcl1d_ca_w_1_360_s_0_360 = 4.53e-05  mcl1d_cc_w_1_360_s_0_360 = 5.82e-11  mcl1d_cf_w_1_360_s_0_360 = 8.35e-12
+ mcl1d_ca_w_1_360_s_0_450 = 4.53e-05  mcl1d_cc_w_1_360_s_0_450 = 5.12e-11  mcl1d_cf_w_1_360_s_0_450 = 1.01e-11
+ mcl1d_ca_w_1_360_s_0_540 = 4.53e-05  mcl1d_cc_w_1_360_s_0_540 = 4.57e-11  mcl1d_cf_w_1_360_s_0_540 = 1.17e-11
+ mcl1d_ca_w_1_360_s_0_720 = 4.53e-05  mcl1d_cc_w_1_360_s_0_720 = 3.80e-11  mcl1d_cf_w_1_360_s_0_720 = 1.48e-11
+ mcl1d_ca_w_1_360_s_1_080 = 4.53e-05  mcl1d_cc_w_1_360_s_1_080 = 2.82e-11  mcl1d_cf_w_1_360_s_1_080 = 1.99e-11
+ mcl1d_ca_w_1_360_s_1_980 = 4.53e-05  mcl1d_cc_w_1_360_s_1_980 = 1.61e-11  mcl1d_cf_w_1_360_s_1_980 = 2.88e-11
+ mcl1d_ca_w_1_360_s_4_500 = 4.53e-05  mcl1d_cc_w_1_360_s_4_500 = 5.75e-12  mcl1d_cf_w_1_360_s_4_500 = 3.82e-11
+ mcl1p1_ca_w_0_170_s_0_180 = 6.45e-05  mcl1p1_cc_w_0_170_s_0_180 = 6.05e-11  mcl1p1_cf_w_0_170_s_0_180 = 6.59e-12
+ mcl1p1_ca_w_0_170_s_0_225 = 6.45e-05  mcl1p1_cc_w_0_170_s_0_225 = 5.24e-11  mcl1p1_cf_w_0_170_s_0_225 = 7.89e-12
+ mcl1p1_ca_w_0_170_s_0_270 = 6.45e-05  mcl1p1_cc_w_0_170_s_0_270 = 4.70e-11  mcl1p1_cf_w_0_170_s_0_270 = 9.11e-12
+ mcl1p1_ca_w_0_170_s_0_360 = 6.45e-05  mcl1p1_cc_w_0_170_s_0_360 = 3.82e-11  mcl1p1_cf_w_0_170_s_0_360 = 1.18e-11
+ mcl1p1_ca_w_0_170_s_0_450 = 6.45e-05  mcl1p1_cc_w_0_170_s_0_450 = 3.28e-11  mcl1p1_cf_w_0_170_s_0_450 = 1.37e-11
+ mcl1p1_ca_w_0_170_s_0_540 = 6.45e-05  mcl1p1_cc_w_0_170_s_0_540 = 2.79e-11  mcl1p1_cf_w_0_170_s_0_540 = 1.60e-11
+ mcl1p1_ca_w_0_170_s_0_720 = 6.45e-05  mcl1p1_cc_w_0_170_s_0_720 = 2.15e-11  mcl1p1_cf_w_0_170_s_0_720 = 1.97e-11
+ mcl1p1_ca_w_0_170_s_1_080 = 6.45e-05  mcl1p1_cc_w_0_170_s_1_080 = 1.40e-11  mcl1p1_cf_w_0_170_s_1_080 = 2.51e-11
+ mcl1p1_ca_w_0_170_s_1_980 = 6.45e-05  mcl1p1_cc_w_0_170_s_1_980 = 6.43e-12  mcl1p1_cf_w_0_170_s_1_980 = 3.16e-11
+ mcl1p1_ca_w_0_170_s_4_500 = 6.45e-05  mcl1p1_cc_w_0_170_s_4_500 = 1.70e-12  mcl1p1_cf_w_0_170_s_4_500 = 3.62e-11
+ mcl1p1_ca_w_1_360_s_0_180 = 6.45e-05  mcl1p1_cc_w_1_360_s_0_180 = 8.01e-11  mcl1p1_cf_w_1_360_s_0_180 = 6.62e-12
+ mcl1p1_ca_w_1_360_s_0_225 = 6.45e-05  mcl1p1_cc_w_1_360_s_0_225 = 7.12e-11  mcl1p1_cf_w_1_360_s_0_225 = 7.92e-12
+ mcl1p1_ca_w_1_360_s_0_270 = 6.45e-05  mcl1p1_cc_w_1_360_s_0_270 = 6.43e-11  mcl1p1_cf_w_1_360_s_0_270 = 9.18e-12
+ mcl1p1_ca_w_1_360_s_0_360 = 6.45e-05  mcl1p1_cc_w_1_360_s_0_360 = 5.42e-11  mcl1p1_cf_w_1_360_s_0_360 = 1.16e-11
+ mcl1p1_ca_w_1_360_s_0_450 = 6.45e-05  mcl1p1_cc_w_1_360_s_0_450 = 4.73e-11  mcl1p1_cf_w_1_360_s_0_450 = 1.39e-11
+ mcl1p1_ca_w_1_360_s_0_540 = 6.45e-05  mcl1p1_cc_w_1_360_s_0_540 = 4.19e-11  mcl1p1_cf_w_1_360_s_0_540 = 1.60e-11
+ mcl1p1_ca_w_1_360_s_0_720 = 6.45e-05  mcl1p1_cc_w_1_360_s_0_720 = 3.42e-11  mcl1p1_cf_w_1_360_s_0_720 = 1.98e-11
+ mcl1p1_ca_w_1_360_s_1_080 = 6.45e-05  mcl1p1_cc_w_1_360_s_1_080 = 2.47e-11  mcl1p1_cf_w_1_360_s_1_080 = 2.59e-11
+ mcl1p1_ca_w_1_360_s_1_980 = 6.45e-05  mcl1p1_cc_w_1_360_s_1_980 = 1.34e-11  mcl1p1_cf_w_1_360_s_1_980 = 3.51e-11
+ mcl1p1_ca_w_1_360_s_4_500 = 6.45e-05  mcl1p1_cc_w_1_360_s_4_500 = 4.55e-12  mcl1p1_cf_w_1_360_s_4_500 = 4.35e-11
+ mcm1f_ca_w_0_140_s_0_140 = 2.02e-05  mcm1f_cc_w_0_140_s_0_140 = 8.80e-11  mcm1f_cf_w_0_140_s_0_140 = 1.70e-12
+ mcm1f_ca_w_0_140_s_0_175 = 2.02e-05  mcm1f_cc_w_0_140_s_0_175 = 8.69e-11  mcm1f_cf_w_0_140_s_0_175 = 2.06e-12
+ mcm1f_ca_w_0_140_s_0_210 = 2.02e-05  mcm1f_cc_w_0_140_s_0_210 = 8.37e-11  mcm1f_cf_w_0_140_s_0_210 = 2.41e-12
+ mcm1f_ca_w_0_140_s_0_280 = 2.02e-05  mcm1f_cc_w_0_140_s_0_280 = 7.60e-11  mcm1f_cf_w_0_140_s_0_280 = 3.10e-12
+ mcm1f_ca_w_0_140_s_0_350 = 2.02e-05  mcm1f_cc_w_0_140_s_0_350 = 6.76e-11  mcm1f_cf_w_0_140_s_0_350 = 3.77e-12
+ mcm1f_ca_w_0_140_s_0_420 = 2.02e-05  mcm1f_cc_w_0_140_s_0_420 = 6.00e-11  mcm1f_cf_w_0_140_s_0_420 = 4.49e-12
+ mcm1f_ca_w_0_140_s_0_560 = 2.02e-05  mcm1f_cc_w_0_140_s_0_560 = 5.05e-11  mcm1f_cf_w_0_140_s_0_560 = 5.75e-12
+ mcm1f_ca_w_0_140_s_0_840 = 2.02e-05  mcm1f_cc_w_0_140_s_0_840 = 3.88e-11  mcm1f_cf_w_0_140_s_0_840 = 8.21e-12
+ mcm1f_ca_w_0_140_s_1_540 = 2.02e-05  mcm1f_cc_w_0_140_s_1_540 = 2.48e-11  mcm1f_cf_w_0_140_s_1_540 = 1.36e-11
+ mcm1f_ca_w_0_140_s_3_500 = 2.02e-05  mcm1f_cc_w_0_140_s_3_500 = 1.09e-11  mcm1f_cf_w_0_140_s_3_500 = 2.29e-11
+ mcm1f_ca_w_1_120_s_0_140 = 2.02e-05  mcm1f_cc_w_1_120_s_0_140 = 1.15e-10  mcm1f_cf_w_1_120_s_0_140 = 1.73e-12
+ mcm1f_ca_w_1_120_s_0_175 = 2.02e-05  mcm1f_cc_w_1_120_s_0_175 = 1.13e-10  mcm1f_cf_w_1_120_s_0_175 = 2.08e-12
+ mcm1f_ca_w_1_120_s_0_210 = 2.02e-05  mcm1f_cc_w_1_120_s_0_210 = 1.08e-10  mcm1f_cf_w_1_120_s_0_210 = 2.43e-12
+ mcm1f_ca_w_1_120_s_0_280 = 2.02e-05  mcm1f_cc_w_1_120_s_0_280 = 9.77e-11  mcm1f_cf_w_1_120_s_0_280 = 3.12e-12
+ mcm1f_ca_w_1_120_s_0_350 = 2.02e-05  mcm1f_cc_w_1_120_s_0_350 = 8.73e-11  mcm1f_cf_w_1_120_s_0_350 = 3.81e-12
+ mcm1f_ca_w_1_120_s_0_420 = 2.02e-05  mcm1f_cc_w_1_120_s_0_420 = 7.84e-11  mcm1f_cf_w_1_120_s_0_420 = 4.48e-12
+ mcm1f_ca_w_1_120_s_0_560 = 2.02e-05  mcm1f_cc_w_1_120_s_0_560 = 6.61e-11  mcm1f_cf_w_1_120_s_0_560 = 5.79e-12
+ mcm1f_ca_w_1_120_s_0_840 = 2.02e-05  mcm1f_cc_w_1_120_s_0_840 = 5.12e-11  mcm1f_cf_w_1_120_s_0_840 = 8.29e-12
+ mcm1f_ca_w_1_120_s_1_540 = 2.02e-05  mcm1f_cc_w_1_120_s_1_540 = 3.37e-11  mcm1f_cf_w_1_120_s_1_540 = 1.39e-11
+ mcm1f_ca_w_1_120_s_3_500 = 2.02e-05  mcm1f_cc_w_1_120_s_3_500 = 1.61e-11  mcm1f_cf_w_1_120_s_3_500 = 2.45e-11
+ mcm1d_ca_w_0_140_s_0_140 = 2.67e-05  mcm1d_cc_w_0_140_s_0_140 = 8.74e-11  mcm1d_cf_w_0_140_s_0_140 = 2.24e-12
+ mcm1d_ca_w_0_140_s_0_175 = 2.67e-05  mcm1d_cc_w_0_140_s_0_175 = 8.60e-11  mcm1d_cf_w_0_140_s_0_175 = 2.71e-12
+ mcm1d_ca_w_0_140_s_0_210 = 2.67e-05  mcm1d_cc_w_0_140_s_0_210 = 8.30e-11  mcm1d_cf_w_0_140_s_0_210 = 3.17e-12
+ mcm1d_ca_w_0_140_s_0_280 = 2.67e-05  mcm1d_cc_w_0_140_s_0_280 = 7.50e-11  mcm1d_cf_w_0_140_s_0_280 = 4.07e-12
+ mcm1d_ca_w_0_140_s_0_350 = 2.67e-05  mcm1d_cc_w_0_140_s_0_350 = 6.63e-11  mcm1d_cf_w_0_140_s_0_350 = 4.94e-12
+ mcm1d_ca_w_0_140_s_0_420 = 2.67e-05  mcm1d_cc_w_0_140_s_0_420 = 5.87e-11  mcm1d_cf_w_0_140_s_0_420 = 5.87e-12
+ mcm1d_ca_w_0_140_s_0_560 = 2.67e-05  mcm1d_cc_w_0_140_s_0_560 = 4.89e-11  mcm1d_cf_w_0_140_s_0_560 = 7.52e-12
+ mcm1d_ca_w_0_140_s_0_840 = 2.67e-05  mcm1d_cc_w_0_140_s_0_840 = 3.68e-11  mcm1d_cf_w_0_140_s_0_840 = 1.06e-11
+ mcm1d_ca_w_0_140_s_1_540 = 2.67e-05  mcm1d_cc_w_0_140_s_1_540 = 2.25e-11  mcm1d_cf_w_0_140_s_1_540 = 1.71e-11
+ mcm1d_ca_w_0_140_s_3_500 = 2.67e-05  mcm1d_cc_w_0_140_s_3_500 = 9.00e-12  mcm1d_cf_w_0_140_s_3_500 = 2.72e-11
+ mcm1d_ca_w_1_120_s_0_140 = 2.67e-05  mcm1d_cc_w_1_120_s_0_140 = 1.13e-10  mcm1d_cf_w_1_120_s_0_140 = 2.28e-12
+ mcm1d_ca_w_1_120_s_0_175 = 2.67e-05  mcm1d_cc_w_1_120_s_0_175 = 1.11e-10  mcm1d_cf_w_1_120_s_0_175 = 2.75e-12
+ mcm1d_ca_w_1_120_s_0_210 = 2.67e-05  mcm1d_cc_w_1_120_s_0_210 = 1.06e-10  mcm1d_cf_w_1_120_s_0_210 = 3.21e-12
+ mcm1d_ca_w_1_120_s_0_280 = 2.67e-05  mcm1d_cc_w_1_120_s_0_280 = 9.51e-11  mcm1d_cf_w_1_120_s_0_280 = 4.11e-12
+ mcm1d_ca_w_1_120_s_0_350 = 2.67e-05  mcm1d_cc_w_1_120_s_0_350 = 8.45e-11  mcm1d_cf_w_1_120_s_0_350 = 5.01e-12
+ mcm1d_ca_w_1_120_s_0_420 = 2.67e-05  mcm1d_cc_w_1_120_s_0_420 = 7.57e-11  mcm1d_cf_w_1_120_s_0_420 = 5.88e-12
+ mcm1d_ca_w_1_120_s_0_560 = 2.67e-05  mcm1d_cc_w_1_120_s_0_560 = 6.34e-11  mcm1d_cf_w_1_120_s_0_560 = 7.57e-12
+ mcm1d_ca_w_1_120_s_0_840 = 2.67e-05  mcm1d_cc_w_1_120_s_0_840 = 4.83e-11  mcm1d_cf_w_1_120_s_0_840 = 1.08e-11
+ mcm1d_ca_w_1_120_s_1_540 = 2.67e-05  mcm1d_cc_w_1_120_s_1_540 = 3.08e-11  mcm1d_cf_w_1_120_s_1_540 = 1.75e-11
+ mcm1d_ca_w_1_120_s_3_500 = 2.67e-05  mcm1d_cc_w_1_120_s_3_500 = 1.37e-11  mcm1d_cf_w_1_120_s_3_500 = 2.93e-11
+ mcm1p1_ca_w_0_140_s_0_140 = 3.23e-05  mcm1p1_cc_w_0_140_s_0_140 = 8.65e-11  mcm1p1_cf_w_0_140_s_0_140 = 2.71e-12
+ mcm1p1_ca_w_0_140_s_0_175 = 3.23e-05  mcm1p1_cc_w_0_140_s_0_175 = 8.53e-11  mcm1p1_cf_w_0_140_s_0_175 = 3.28e-12
+ mcm1p1_ca_w_0_140_s_0_210 = 3.23e-05  mcm1p1_cc_w_0_140_s_0_210 = 8.22e-11  mcm1p1_cf_w_0_140_s_0_210 = 3.83e-12
+ mcm1p1_ca_w_0_140_s_0_280 = 3.23e-05  mcm1p1_cc_w_0_140_s_0_280 = 7.41e-11  mcm1p1_cf_w_0_140_s_0_280 = 4.93e-12
+ mcm1p1_ca_w_0_140_s_0_350 = 3.23e-05  mcm1p1_cc_w_0_140_s_0_350 = 6.51e-11  mcm1p1_cf_w_0_140_s_0_350 = 5.98e-12
+ mcm1p1_ca_w_0_140_s_0_420 = 3.23e-05  mcm1p1_cc_w_0_140_s_0_420 = 5.78e-11  mcm1p1_cf_w_0_140_s_0_420 = 7.06e-12
+ mcm1p1_ca_w_0_140_s_0_560 = 3.23e-05  mcm1p1_cc_w_0_140_s_0_560 = 4.75e-11  mcm1p1_cf_w_0_140_s_0_560 = 9.02e-12
+ mcm1p1_ca_w_0_140_s_0_840 = 3.23e-05  mcm1p1_cc_w_0_140_s_0_840 = 3.52e-11  mcm1p1_cf_w_0_140_s_0_840 = 1.27e-11
+ mcm1p1_ca_w_0_140_s_1_540 = 3.23e-05  mcm1p1_cc_w_0_140_s_1_540 = 2.07e-11  mcm1p1_cf_w_0_140_s_1_540 = 2.00e-11
+ mcm1p1_ca_w_0_140_s_3_500 = 3.23e-05  mcm1p1_cc_w_0_140_s_3_500 = 7.74e-12  mcm1p1_cf_w_0_140_s_3_500 = 3.03e-11
+ mcm1p1_ca_w_1_120_s_0_140 = 3.23e-05  mcm1p1_cc_w_1_120_s_0_140 = 1.11e-10  mcm1p1_cf_w_1_120_s_0_140 = 2.80e-12
+ mcm1p1_ca_w_1_120_s_0_175 = 3.23e-05  mcm1p1_cc_w_1_120_s_0_175 = 1.08e-10  mcm1p1_cf_w_1_120_s_0_175 = 3.36e-12
+ mcm1p1_ca_w_1_120_s_0_210 = 3.23e-05  mcm1p1_cc_w_1_120_s_0_210 = 1.04e-10  mcm1p1_cf_w_1_120_s_0_210 = 3.90e-12
+ mcm1p1_ca_w_1_120_s_0_280 = 3.23e-05  mcm1p1_cc_w_1_120_s_0_280 = 9.30e-11  mcm1p1_cf_w_1_120_s_0_280 = 5.01e-12
+ mcm1p1_ca_w_1_120_s_0_350 = 3.23e-05  mcm1p1_cc_w_1_120_s_0_350 = 8.28e-11  mcm1p1_cf_w_1_120_s_0_350 = 6.08e-12
+ mcm1p1_ca_w_1_120_s_0_420 = 3.23e-05  mcm1p1_cc_w_1_120_s_0_420 = 7.39e-11  mcm1p1_cf_w_1_120_s_0_420 = 7.12e-12
+ mcm1p1_ca_w_1_120_s_0_560 = 3.23e-05  mcm1p1_cc_w_1_120_s_0_560 = 6.12e-11  mcm1p1_cf_w_1_120_s_0_560 = 9.12e-12
+ mcm1p1_ca_w_1_120_s_0_840 = 3.23e-05  mcm1p1_cc_w_1_120_s_0_840 = 4.62e-11  mcm1p1_cf_w_1_120_s_0_840 = 1.28e-11
+ mcm1p1_ca_w_1_120_s_1_540 = 3.23e-05  mcm1p1_cc_w_1_120_s_1_540 = 2.87e-11  mcm1p1_cf_w_1_120_s_1_540 = 2.06e-11
+ mcm1p1_ca_w_1_120_s_3_500 = 3.23e-05  mcm1p1_cc_w_1_120_s_3_500 = 1.22e-11  mcm1p1_cf_w_1_120_s_3_500 = 3.28e-11
+ mcm1l1_ca_w_0_140_s_0_140 = 7.72e-05  mcm1l1_cc_w_0_140_s_0_140 = 8.19e-11  mcm1l1_cf_w_0_140_s_0_140 = 6.21e-12
+ mcm1l1_ca_w_0_140_s_0_175 = 7.72e-05  mcm1l1_cc_w_0_140_s_0_175 = 8.04e-11  mcm1l1_cf_w_0_140_s_0_175 = 7.56e-12
+ mcm1l1_ca_w_0_140_s_0_210 = 7.72e-05  mcm1l1_cc_w_0_140_s_0_210 = 7.71e-11  mcm1l1_cf_w_0_140_s_0_210 = 8.84e-12
+ mcm1l1_ca_w_0_140_s_0_280 = 7.72e-05  mcm1l1_cc_w_0_140_s_0_280 = 6.81e-11  mcm1l1_cf_w_0_140_s_0_280 = 1.13e-11
+ mcm1l1_ca_w_0_140_s_0_350 = 7.72e-05  mcm1l1_cc_w_0_140_s_0_350 = 5.86e-11  mcm1l1_cf_w_0_140_s_0_350 = 1.36e-11
+ mcm1l1_ca_w_0_140_s_0_420 = 7.72e-05  mcm1l1_cc_w_0_140_s_0_420 = 5.07e-11  mcm1l1_cf_w_0_140_s_0_420 = 1.59e-11
+ mcm1l1_ca_w_0_140_s_0_560 = 7.72e-05  mcm1l1_cc_w_0_140_s_0_560 = 3.99e-11  mcm1l1_cf_w_0_140_s_0_560 = 1.99e-11
+ mcm1l1_ca_w_0_140_s_0_840 = 7.72e-05  mcm1l1_cc_w_0_140_s_0_840 = 2.72e-11  mcm1l1_cf_w_0_140_s_0_840 = 2.64e-11
+ mcm1l1_ca_w_0_140_s_1_540 = 7.72e-05  mcm1l1_cc_w_0_140_s_1_540 = 1.35e-11  mcm1l1_cf_w_0_140_s_1_540 = 3.68e-11
+ mcm1l1_ca_w_0_140_s_3_500 = 7.72e-05  mcm1l1_cc_w_0_140_s_3_500 = 3.97e-12  mcm1l1_cf_w_0_140_s_3_500 = 4.58e-11
+ mcm1l1_ca_w_1_120_s_0_140 = 7.72e-05  mcm1l1_cc_w_1_120_s_0_140 = 1.01e-10  mcm1l1_cf_w_1_120_s_0_140 = 6.29e-12
+ mcm1l1_ca_w_1_120_s_0_175 = 7.72e-05  mcm1l1_cc_w_1_120_s_0_175 = 9.86e-11  mcm1l1_cf_w_1_120_s_0_175 = 7.62e-12
+ mcm1l1_ca_w_1_120_s_0_210 = 7.72e-05  mcm1l1_cc_w_1_120_s_0_210 = 9.39e-11  mcm1l1_cf_w_1_120_s_0_210 = 8.92e-12
+ mcm1l1_ca_w_1_120_s_0_280 = 7.72e-05  mcm1l1_cc_w_1_120_s_0_280 = 8.30e-11  mcm1l1_cf_w_1_120_s_0_280 = 1.14e-11
+ mcm1l1_ca_w_1_120_s_0_350 = 7.72e-05  mcm1l1_cc_w_1_120_s_0_350 = 7.31e-11  mcm1l1_cf_w_1_120_s_0_350 = 1.37e-11
+ mcm1l1_ca_w_1_120_s_0_420 = 7.72e-05  mcm1l1_cc_w_1_120_s_0_420 = 6.40e-11  mcm1l1_cf_w_1_120_s_0_420 = 1.59e-11
+ mcm1l1_ca_w_1_120_s_0_560 = 7.72e-05  mcm1l1_cc_w_1_120_s_0_560 = 5.16e-11  mcm1l1_cf_w_1_120_s_0_560 = 1.99e-11
+ mcm1l1_ca_w_1_120_s_0_840 = 7.72e-05  mcm1l1_cc_w_1_120_s_0_840 = 3.71e-11  mcm1l1_cf_w_1_120_s_0_840 = 2.67e-11
+ mcm1l1_ca_w_1_120_s_1_540 = 7.72e-05  mcm1l1_cc_w_1_120_s_1_540 = 2.08e-11  mcm1l1_cf_w_1_120_s_1_540 = 3.77e-11
+ mcm1l1_ca_w_1_120_s_3_500 = 7.72e-05  mcm1l1_cc_w_1_120_s_3_500 = 7.60e-12  mcm1l1_cf_w_1_120_s_3_500 = 4.97e-11
+ mcm2f_ca_w_0_140_s_0_140 = 1.40e-05  mcm2f_cc_w_0_140_s_0_140 = 8.86e-11  mcm2f_cf_w_0_140_s_0_140 = 1.19e-12
+ mcm2f_ca_w_0_140_s_0_175 = 1.40e-05  mcm2f_cc_w_0_140_s_0_175 = 8.74e-11  mcm2f_cf_w_0_140_s_0_175 = 1.43e-12
+ mcm2f_ca_w_0_140_s_0_210 = 1.40e-05  mcm2f_cc_w_0_140_s_0_210 = 8.46e-11  mcm2f_cf_w_0_140_s_0_210 = 1.68e-12
+ mcm2f_ca_w_0_140_s_0_280 = 1.40e-05  mcm2f_cc_w_0_140_s_0_280 = 7.71e-11  mcm2f_cf_w_0_140_s_0_280 = 2.16e-12
+ mcm2f_ca_w_0_140_s_0_350 = 1.40e-05  mcm2f_cc_w_0_140_s_0_350 = 6.86e-11  mcm2f_cf_w_0_140_s_0_350 = 2.63e-12
+ mcm2f_ca_w_0_140_s_0_420 = 1.40e-05  mcm2f_cc_w_0_140_s_0_420 = 6.13e-11  mcm2f_cf_w_0_140_s_0_420 = 3.13e-12
+ mcm2f_ca_w_0_140_s_0_560 = 1.40e-05  mcm2f_cc_w_0_140_s_0_560 = 5.18e-11  mcm2f_cf_w_0_140_s_0_560 = 4.02e-12
+ mcm2f_ca_w_0_140_s_0_840 = 1.40e-05  mcm2f_cc_w_0_140_s_0_840 = 4.06e-11  mcm2f_cf_w_0_140_s_0_840 = 5.80e-12
+ mcm2f_ca_w_0_140_s_1_540 = 1.40e-05  mcm2f_cc_w_0_140_s_1_540 = 2.73e-11  mcm2f_cf_w_0_140_s_1_540 = 9.83e-12
+ mcm2f_ca_w_0_140_s_3_500 = 1.40e-05  mcm2f_cc_w_0_140_s_3_500 = 1.36e-11  mcm2f_cf_w_0_140_s_3_500 = 1.78e-11
+ mcm2f_ca_w_1_120_s_0_140 = 1.40e-05  mcm2f_cc_w_1_120_s_0_140 = 1.18e-10  mcm2f_cf_w_1_120_s_0_140 = 1.20e-12
+ mcm2f_ca_w_1_120_s_0_175 = 1.40e-05  mcm2f_cc_w_1_120_s_0_175 = 1.15e-10  mcm2f_cf_w_1_120_s_0_175 = 1.45e-12
+ mcm2f_ca_w_1_120_s_0_210 = 1.40e-05  mcm2f_cc_w_1_120_s_0_210 = 1.11e-10  mcm2f_cf_w_1_120_s_0_210 = 1.69e-12
+ mcm2f_ca_w_1_120_s_0_280 = 1.40e-05  mcm2f_cc_w_1_120_s_0_280 = 9.97e-11  mcm2f_cf_w_1_120_s_0_280 = 2.17e-12
+ mcm2f_ca_w_1_120_s_0_350 = 1.40e-05  mcm2f_cc_w_1_120_s_0_350 = 8.98e-11  mcm2f_cf_w_1_120_s_0_350 = 2.65e-12
+ mcm2f_ca_w_1_120_s_0_420 = 1.40e-05  mcm2f_cc_w_1_120_s_0_420 = 8.09e-11  mcm2f_cf_w_1_120_s_0_420 = 3.12e-12
+ mcm2f_ca_w_1_120_s_0_560 = 1.40e-05  mcm2f_cc_w_1_120_s_0_560 = 6.87e-11  mcm2f_cf_w_1_120_s_0_560 = 4.05e-12
+ mcm2f_ca_w_1_120_s_0_840 = 1.40e-05  mcm2f_cc_w_1_120_s_0_840 = 5.41e-11  mcm2f_cf_w_1_120_s_0_840 = 5.86e-12
+ mcm2f_ca_w_1_120_s_1_540 = 1.40e-05  mcm2f_cc_w_1_120_s_1_540 = 3.68e-11  mcm2f_cf_w_1_120_s_1_540 = 9.99e-12
+ mcm2f_ca_w_1_120_s_3_500 = 1.40e-05  mcm2f_cc_w_1_120_s_3_500 = 1.93e-11  mcm2f_cf_w_1_120_s_3_500 = 1.89e-11
+ mcm2d_ca_w_0_140_s_0_140 = 1.68e-05  mcm2d_cc_w_0_140_s_0_140 = 8.84e-11  mcm2d_cf_w_0_140_s_0_140 = 1.42e-12
+ mcm2d_ca_w_0_140_s_0_175 = 1.68e-05  mcm2d_cc_w_0_140_s_0_175 = 8.70e-11  mcm2d_cf_w_0_140_s_0_175 = 1.71e-12
+ mcm2d_ca_w_0_140_s_0_210 = 1.68e-05  mcm2d_cc_w_0_140_s_0_210 = 8.42e-11  mcm2d_cf_w_0_140_s_0_210 = 2.01e-12
+ mcm2d_ca_w_0_140_s_0_280 = 1.68e-05  mcm2d_cc_w_0_140_s_0_280 = 7.66e-11  mcm2d_cf_w_0_140_s_0_280 = 2.59e-12
+ mcm2d_ca_w_0_140_s_0_350 = 1.68e-05  mcm2d_cc_w_0_140_s_0_350 = 6.79e-11  mcm2d_cf_w_0_140_s_0_350 = 3.15e-12
+ mcm2d_ca_w_0_140_s_0_420 = 1.68e-05  mcm2d_cc_w_0_140_s_0_420 = 6.06e-11  mcm2d_cf_w_0_140_s_0_420 = 3.74e-12
+ mcm2d_ca_w_0_140_s_0_560 = 1.68e-05  mcm2d_cc_w_0_140_s_0_560 = 5.10e-11  mcm2d_cf_w_0_140_s_0_560 = 4.80e-12
+ mcm2d_ca_w_0_140_s_0_840 = 1.68e-05  mcm2d_cc_w_0_140_s_0_840 = 3.96e-11  mcm2d_cf_w_0_140_s_0_840 = 6.91e-12
+ mcm2d_ca_w_0_140_s_1_540 = 1.68e-05  mcm2d_cc_w_0_140_s_1_540 = 2.60e-11  mcm2d_cf_w_0_140_s_1_540 = 1.16e-11
+ mcm2d_ca_w_0_140_s_3_500 = 1.68e-05  mcm2d_cc_w_0_140_s_3_500 = 1.22e-11  mcm2d_cf_w_0_140_s_3_500 = 2.03e-11
+ mcm2d_ca_w_1_120_s_0_140 = 1.68e-05  mcm2d_cc_w_1_120_s_0_140 = 1.16e-10  mcm2d_cf_w_1_120_s_0_140 = 1.45e-12
+ mcm2d_ca_w_1_120_s_0_175 = 1.68e-05  mcm2d_cc_w_1_120_s_0_175 = 1.14e-10  mcm2d_cf_w_1_120_s_0_175 = 1.74e-12
+ mcm2d_ca_w_1_120_s_0_210 = 1.68e-05  mcm2d_cc_w_1_120_s_0_210 = 1.10e-10  mcm2d_cf_w_1_120_s_0_210 = 2.03e-12
+ mcm2d_ca_w_1_120_s_0_280 = 1.68e-05  mcm2d_cc_w_1_120_s_0_280 = 9.83e-11  mcm2d_cf_w_1_120_s_0_280 = 2.61e-12
+ mcm2d_ca_w_1_120_s_0_350 = 1.68e-05  mcm2d_cc_w_1_120_s_0_350 = 8.84e-11  mcm2d_cf_w_1_120_s_0_350 = 3.18e-12
+ mcm2d_ca_w_1_120_s_0_420 = 1.68e-05  mcm2d_cc_w_1_120_s_0_420 = 7.94e-11  mcm2d_cf_w_1_120_s_0_420 = 3.75e-12
+ mcm2d_ca_w_1_120_s_0_560 = 1.68e-05  mcm2d_cc_w_1_120_s_0_560 = 6.72e-11  mcm2d_cf_w_1_120_s_0_560 = 4.85e-12
+ mcm2d_ca_w_1_120_s_0_840 = 1.68e-05  mcm2d_cc_w_1_120_s_0_840 = 5.24e-11  mcm2d_cf_w_1_120_s_0_840 = 6.98e-12
+ mcm2d_ca_w_1_120_s_1_540 = 1.68e-05  mcm2d_cc_w_1_120_s_1_540 = 3.51e-11  mcm2d_cf_w_1_120_s_1_540 = 1.18e-11
+ mcm2d_ca_w_1_120_s_3_500 = 1.68e-05  mcm2d_cc_w_1_120_s_3_500 = 1.75e-11  mcm2d_cf_w_1_120_s_3_500 = 2.16e-11
+ mcm2p1_ca_w_0_140_s_0_140 = 1.89e-05  mcm2p1_cc_w_0_140_s_0_140 = 8.79e-11  mcm2p1_cf_w_0_140_s_0_140 = 1.60e-12
+ mcm2p1_ca_w_0_140_s_0_175 = 1.89e-05  mcm2p1_cc_w_0_140_s_0_175 = 8.67e-11  mcm2p1_cf_w_0_140_s_0_175 = 1.93e-12
+ mcm2p1_ca_w_0_140_s_0_210 = 1.89e-05  mcm2p1_cc_w_0_140_s_0_210 = 8.39e-11  mcm2p1_cf_w_0_140_s_0_210 = 2.26e-12
+ mcm2p1_ca_w_0_140_s_0_280 = 1.89e-05  mcm2p1_cc_w_0_140_s_0_280 = 7.62e-11  mcm2p1_cf_w_0_140_s_0_280 = 2.91e-12
+ mcm2p1_ca_w_0_140_s_0_350 = 1.89e-05  mcm2p1_cc_w_0_140_s_0_350 = 6.75e-11  mcm2p1_cf_w_0_140_s_0_350 = 3.54e-12
+ mcm2p1_ca_w_0_140_s_0_420 = 1.89e-05  mcm2p1_cc_w_0_140_s_0_420 = 6.05e-11  mcm2p1_cf_w_0_140_s_0_420 = 4.20e-12
+ mcm2p1_ca_w_0_140_s_0_560 = 1.89e-05  mcm2p1_cc_w_0_140_s_0_560 = 5.05e-11  mcm2p1_cf_w_0_140_s_0_560 = 5.39e-12
+ mcm2p1_ca_w_0_140_s_0_840 = 1.89e-05  mcm2p1_cc_w_0_140_s_0_840 = 3.89e-11  mcm2p1_cf_w_0_140_s_0_840 = 7.73e-12
+ mcm2p1_ca_w_0_140_s_1_540 = 1.89e-05  mcm2p1_cc_w_0_140_s_1_540 = 2.51e-11  mcm2p1_cf_w_0_140_s_1_540 = 1.28e-11
+ mcm2p1_ca_w_0_140_s_3_500 = 1.89e-05  mcm2p1_cc_w_0_140_s_3_500 = 1.13e-11  mcm2p1_cf_w_0_140_s_3_500 = 2.19e-11
+ mcm2p1_ca_w_1_120_s_0_140 = 1.89e-05  mcm2p1_cc_w_1_120_s_0_140 = 1.16e-10  mcm2p1_cf_w_1_120_s_0_140 = 1.64e-12
+ mcm2p1_ca_w_1_120_s_0_175 = 1.89e-05  mcm2p1_cc_w_1_120_s_0_175 = 1.13e-10  mcm2p1_cf_w_1_120_s_0_175 = 1.97e-12
+ mcm2p1_ca_w_1_120_s_0_210 = 1.89e-05  mcm2p1_cc_w_1_120_s_0_210 = 1.09e-10  mcm2p1_cf_w_1_120_s_0_210 = 2.30e-12
+ mcm2p1_ca_w_1_120_s_0_280 = 1.89e-05  mcm2p1_cc_w_1_120_s_0_280 = 9.73e-11  mcm2p1_cf_w_1_120_s_0_280 = 2.95e-12
+ mcm2p1_ca_w_1_120_s_0_350 = 1.89e-05  mcm2p1_cc_w_1_120_s_0_350 = 8.74e-11  mcm2p1_cf_w_1_120_s_0_350 = 3.59e-12
+ mcm2p1_ca_w_1_120_s_0_420 = 1.89e-05  mcm2p1_cc_w_1_120_s_0_420 = 7.87e-11  mcm2p1_cf_w_1_120_s_0_420 = 4.23e-12
+ mcm2p1_ca_w_1_120_s_0_560 = 1.89e-05  mcm2p1_cc_w_1_120_s_0_560 = 6.62e-11  mcm2p1_cf_w_1_120_s_0_560 = 5.45e-12
+ mcm2p1_ca_w_1_120_s_0_840 = 1.89e-05  mcm2p1_cc_w_1_120_s_0_840 = 5.13e-11  mcm2p1_cf_w_1_120_s_0_840 = 7.82e-12
+ mcm2p1_ca_w_1_120_s_1_540 = 1.89e-05  mcm2p1_cc_w_1_120_s_1_540 = 3.39e-11  mcm2p1_cf_w_1_120_s_1_540 = 1.31e-11
+ mcm2p1_ca_w_1_120_s_3_500 = 1.89e-05  mcm2p1_cc_w_1_120_s_3_500 = 1.64e-11  mcm2p1_cf_w_1_120_s_3_500 = 2.34e-11
+ mcm2l1_ca_w_0_140_s_0_140 = 2.86e-05  mcm2l1_cc_w_0_140_s_0_140 = 8.68e-11  mcm2l1_cf_w_0_140_s_0_140 = 2.40e-12
+ mcm2l1_ca_w_0_140_s_0_175 = 2.86e-05  mcm2l1_cc_w_0_140_s_0_175 = 8.57e-11  mcm2l1_cf_w_0_140_s_0_175 = 2.90e-12
+ mcm2l1_ca_w_0_140_s_0_210 = 2.86e-05  mcm2l1_cc_w_0_140_s_0_210 = 8.27e-11  mcm2l1_cf_w_0_140_s_0_210 = 3.39e-12
+ mcm2l1_ca_w_0_140_s_0_280 = 2.86e-05  mcm2l1_cc_w_0_140_s_0_280 = 7.46e-11  mcm2l1_cf_w_0_140_s_0_280 = 4.36e-12
+ mcm2l1_ca_w_0_140_s_0_350 = 2.86e-05  mcm2l1_cc_w_0_140_s_0_350 = 6.57e-11  mcm2l1_cf_w_0_140_s_0_350 = 5.29e-12
+ mcm2l1_ca_w_0_140_s_0_420 = 2.86e-05  mcm2l1_cc_w_0_140_s_0_420 = 5.85e-11  mcm2l1_cf_w_0_140_s_0_420 = 6.25e-12
+ mcm2l1_ca_w_0_140_s_0_560 = 2.86e-05  mcm2l1_cc_w_0_140_s_0_560 = 4.82e-11  mcm2l1_cf_w_0_140_s_0_560 = 8.01e-12
+ mcm2l1_ca_w_0_140_s_0_840 = 2.86e-05  mcm2l1_cc_w_0_140_s_0_840 = 3.60e-11  mcm2l1_cf_w_0_140_s_0_840 = 1.13e-11
+ mcm2l1_ca_w_0_140_s_1_540 = 2.86e-05  mcm2l1_cc_w_0_140_s_1_540 = 2.16e-11  mcm2l1_cf_w_0_140_s_1_540 = 1.81e-11
+ mcm2l1_ca_w_0_140_s_3_500 = 2.86e-05  mcm2l1_cc_w_0_140_s_3_500 = 8.41e-12  mcm2l1_cf_w_0_140_s_3_500 = 2.82e-11
+ mcm2l1_ca_w_1_120_s_0_140 = 2.86e-05  mcm2l1_cc_w_1_120_s_0_140 = 1.12e-10  mcm2l1_cf_w_1_120_s_0_140 = 2.42e-12
+ mcm2l1_ca_w_1_120_s_0_175 = 2.86e-05  mcm2l1_cc_w_1_120_s_0_175 = 1.09e-10  mcm2l1_cf_w_1_120_s_0_175 = 2.92e-12
+ mcm2l1_ca_w_1_120_s_0_210 = 2.86e-05  mcm2l1_cc_w_1_120_s_0_210 = 1.05e-10  mcm2l1_cf_w_1_120_s_0_210 = 3.41e-12
+ mcm2l1_ca_w_1_120_s_0_280 = 2.86e-05  mcm2l1_cc_w_1_120_s_0_280 = 9.40e-11  mcm2l1_cf_w_1_120_s_0_280 = 4.38e-12
+ mcm2l1_ca_w_1_120_s_0_350 = 2.86e-05  mcm2l1_cc_w_1_120_s_0_350 = 8.35e-11  mcm2l1_cf_w_1_120_s_0_350 = 5.34e-12
+ mcm2l1_ca_w_1_120_s_0_420 = 2.86e-05  mcm2l1_cc_w_1_120_s_0_420 = 7.48e-11  mcm2l1_cf_w_1_120_s_0_420 = 6.26e-12
+ mcm2l1_ca_w_1_120_s_0_560 = 2.86e-05  mcm2l1_cc_w_1_120_s_0_560 = 6.21e-11  mcm2l1_cf_w_1_120_s_0_560 = 8.07e-12
+ mcm2l1_ca_w_1_120_s_0_840 = 2.86e-05  mcm2l1_cc_w_1_120_s_0_840 = 4.72e-11  mcm2l1_cf_w_1_120_s_0_840 = 1.14e-11
+ mcm2l1_ca_w_1_120_s_1_540 = 2.86e-05  mcm2l1_cc_w_1_120_s_1_540 = 2.96e-11  mcm2l1_cf_w_1_120_s_1_540 = 1.85e-11
+ mcm2l1_ca_w_1_120_s_3_500 = 2.86e-05  mcm2l1_cc_w_1_120_s_3_500 = 1.30e-11  mcm2l1_cf_w_1_120_s_3_500 = 3.03e-11
+ mcm2m1_ca_w_0_140_s_0_140 = 8.04e-05  mcm2m1_cc_w_0_140_s_0_140 = 8.14e-11  mcm2m1_cf_w_0_140_s_0_140 = 6.42e-12
+ mcm2m1_ca_w_0_140_s_0_175 = 8.04e-05  mcm2m1_cc_w_0_140_s_0_175 = 8.01e-11  mcm2m1_cf_w_0_140_s_0_175 = 7.82e-12
+ mcm2m1_ca_w_0_140_s_0_210 = 8.04e-05  mcm2m1_cc_w_0_140_s_0_210 = 7.68e-11  mcm2m1_cf_w_0_140_s_0_210 = 9.16e-12
+ mcm2m1_ca_w_0_140_s_0_280 = 8.04e-05  mcm2m1_cc_w_0_140_s_0_280 = 6.78e-11  mcm2m1_cf_w_0_140_s_0_280 = 1.17e-11
+ mcm2m1_ca_w_0_140_s_0_350 = 8.04e-05  mcm2m1_cc_w_0_140_s_0_350 = 5.83e-11  mcm2m1_cf_w_0_140_s_0_350 = 1.41e-11
+ mcm2m1_ca_w_0_140_s_0_420 = 8.04e-05  mcm2m1_cc_w_0_140_s_0_420 = 5.03e-11  mcm2m1_cf_w_0_140_s_0_420 = 1.64e-11
+ mcm2m1_ca_w_0_140_s_0_560 = 8.04e-05  mcm2m1_cc_w_0_140_s_0_560 = 3.95e-11  mcm2m1_cf_w_0_140_s_0_560 = 2.05e-11
+ mcm2m1_ca_w_0_140_s_0_840 = 8.04e-05  mcm2m1_cc_w_0_140_s_0_840 = 2.69e-11  mcm2m1_cf_w_0_140_s_0_840 = 2.72e-11
+ mcm2m1_ca_w_0_140_s_1_540 = 8.04e-05  mcm2m1_cc_w_0_140_s_1_540 = 1.32e-11  mcm2m1_cf_w_0_140_s_1_540 = 3.77e-11
+ mcm2m1_ca_w_0_140_s_3_500 = 8.04e-05  mcm2m1_cc_w_0_140_s_3_500 = 3.85e-12  mcm2m1_cf_w_0_140_s_3_500 = 4.65e-11
+ mcm2m1_ca_w_1_120_s_0_140 = 8.04e-05  mcm2m1_cc_w_1_120_s_0_140 = 1.01e-10  mcm2m1_cf_w_1_120_s_0_140 = 6.45e-12
+ mcm2m1_ca_w_1_120_s_0_175 = 8.04e-05  mcm2m1_cc_w_1_120_s_0_175 = 9.81e-11  mcm2m1_cf_w_1_120_s_0_175 = 7.84e-12
+ mcm2m1_ca_w_1_120_s_0_210 = 8.04e-05  mcm2m1_cc_w_1_120_s_0_210 = 9.35e-11  mcm2m1_cf_w_1_120_s_0_210 = 9.18e-12
+ mcm2m1_ca_w_1_120_s_0_280 = 8.04e-05  mcm2m1_cc_w_1_120_s_0_280 = 8.27e-11  mcm2m1_cf_w_1_120_s_0_280 = 1.17e-11
+ mcm2m1_ca_w_1_120_s_0_350 = 8.04e-05  mcm2m1_cc_w_1_120_s_0_350 = 7.23e-11  mcm2m1_cf_w_1_120_s_0_350 = 1.41e-11
+ mcm2m1_ca_w_1_120_s_0_420 = 8.04e-05  mcm2m1_cc_w_1_120_s_0_420 = 6.36e-11  mcm2m1_cf_w_1_120_s_0_420 = 1.64e-11
+ mcm2m1_ca_w_1_120_s_0_560 = 8.04e-05  mcm2m1_cc_w_1_120_s_0_560 = 5.13e-11  mcm2m1_cf_w_1_120_s_0_560 = 2.06e-11
+ mcm2m1_ca_w_1_120_s_0_840 = 8.04e-05  mcm2m1_cc_w_1_120_s_0_840 = 3.68e-11  mcm2m1_cf_w_1_120_s_0_840 = 2.74e-11
+ mcm2m1_ca_w_1_120_s_1_540 = 8.04e-05  mcm2m1_cc_w_1_120_s_1_540 = 2.05e-11  mcm2m1_cf_w_1_120_s_1_540 = 3.86e-11
+ mcm2m1_ca_w_1_120_s_3_500 = 8.04e-05  mcm2m1_cc_w_1_120_s_3_500 = 7.50e-12  mcm2m1_cf_w_1_120_s_3_500 = 5.04e-11
+ mcm3f_ca_w_0_300_s_0_300 = 1.02e-05  mcm3f_cc_w_0_300_s_0_300 = 9.20e-11  mcm3f_cf_w_0_300_s_0_300 = 1.75e-12
+ mcm3f_ca_w_0_300_s_0_360 = 1.02e-05  mcm3f_cc_w_0_300_s_0_360 = 8.67e-11  mcm3f_cf_w_0_300_s_0_360 = 2.05e-12
+ mcm3f_ca_w_0_300_s_0_450 = 1.02e-05  mcm3f_cc_w_0_300_s_0_450 = 7.91e-11  mcm3f_cf_w_0_300_s_0_450 = 2.52e-12
+ mcm3f_ca_w_0_300_s_0_600 = 1.02e-05  mcm3f_cc_w_0_300_s_0_600 = 6.91e-11  mcm3f_cf_w_0_300_s_0_600 = 3.27e-12
+ mcm3f_ca_w_0_300_s_0_800 = 1.02e-05  mcm3f_cc_w_0_300_s_0_800 = 5.94e-11  mcm3f_cf_w_0_300_s_0_800 = 4.15e-12
+ mcm3f_ca_w_0_300_s_1_000 = 1.02e-05  mcm3f_cc_w_0_300_s_1_000 = 5.20e-11  mcm3f_cf_w_0_300_s_1_000 = 5.08e-12
+ mcm3f_ca_w_0_300_s_1_200 = 1.02e-05  mcm3f_cc_w_0_300_s_1_200 = 4.63e-11  mcm3f_cf_w_0_300_s_1_200 = 5.97e-12
+ mcm3f_ca_w_0_300_s_2_100 = 1.02e-05  mcm3f_cc_w_0_300_s_2_100 = 3.15e-11  mcm3f_cf_w_0_300_s_2_100 = 1.00e-11
+ mcm3f_ca_w_0_300_s_3_300 = 1.02e-05  mcm3f_cc_w_0_300_s_3_300 = 2.25e-11  mcm3f_cf_w_0_300_s_3_300 = 1.39e-11
+ mcm3f_ca_w_0_300_s_9_000 = 1.02e-05  mcm3f_cc_w_0_300_s_9_000 = 7.39e-12  mcm3f_cf_w_0_300_s_9_000 = 2.48e-11
+ mcm3f_ca_w_2_400_s_0_300 = 1.02e-05  mcm3f_cc_w_2_400_s_0_300 = 1.18e-10  mcm3f_cf_w_2_400_s_0_300 = 1.78e-12
+ mcm3f_ca_w_2_400_s_0_360 = 1.02e-05  mcm3f_cc_w_2_400_s_0_360 = 1.12e-10  mcm3f_cf_w_2_400_s_0_360 = 2.07e-12
+ mcm3f_ca_w_2_400_s_0_450 = 1.02e-05  mcm3f_cc_w_2_400_s_0_450 = 1.03e-10  mcm3f_cf_w_2_400_s_0_450 = 2.52e-12
+ mcm3f_ca_w_2_400_s_0_600 = 1.02e-05  mcm3f_cc_w_2_400_s_0_600 = 9.05e-11  mcm3f_cf_w_2_400_s_0_600 = 3.25e-12
+ mcm3f_ca_w_2_400_s_0_800 = 1.02e-05  mcm3f_cc_w_2_400_s_0_800 = 7.82e-11  mcm3f_cf_w_2_400_s_0_800 = 4.20e-12
+ mcm3f_ca_w_2_400_s_1_000 = 1.02e-05  mcm3f_cc_w_2_400_s_1_000 = 6.87e-11  mcm3f_cf_w_2_400_s_1_000 = 5.14e-12
+ mcm3f_ca_w_2_400_s_1_200 = 1.02e-05  mcm3f_cc_w_2_400_s_1_200 = 6.16e-11  mcm3f_cf_w_2_400_s_1_200 = 6.05e-12
+ mcm3f_ca_w_2_400_s_2_100 = 1.02e-05  mcm3f_cc_w_2_400_s_2_100 = 4.32e-11  mcm3f_cf_w_2_400_s_2_100 = 9.91e-12
+ mcm3f_ca_w_2_400_s_3_300 = 1.02e-05  mcm3f_cc_w_2_400_s_3_300 = 3.12e-11  mcm3f_cf_w_2_400_s_3_300 = 1.44e-11
+ mcm3f_ca_w_2_400_s_9_000 = 1.02e-05  mcm3f_cc_w_2_400_s_9_000 = 1.14e-11  mcm3f_cf_w_2_400_s_9_000 = 2.74e-11
+ mcm3d_ca_w_0_300_s_0_300 = 1.17e-05  mcm3d_cc_w_0_300_s_0_300 = 9.15e-11  mcm3d_cf_w_0_300_s_0_300 = 1.99e-12
+ mcm3d_ca_w_0_300_s_0_360 = 1.17e-05  mcm3d_cc_w_0_300_s_0_360 = 8.63e-11  mcm3d_cf_w_0_300_s_0_360 = 2.33e-12
+ mcm3d_ca_w_0_300_s_0_450 = 1.17e-05  mcm3d_cc_w_0_300_s_0_450 = 7.87e-11  mcm3d_cf_w_0_300_s_0_450 = 2.86e-12
+ mcm3d_ca_w_0_300_s_0_600 = 1.17e-05  mcm3d_cc_w_0_300_s_0_600 = 6.86e-11  mcm3d_cf_w_0_300_s_0_600 = 3.71e-12
+ mcm3d_ca_w_0_300_s_0_800 = 1.17e-05  mcm3d_cc_w_0_300_s_0_800 = 5.88e-11  mcm3d_cf_w_0_300_s_0_800 = 4.71e-12
+ mcm3d_ca_w_0_300_s_1_000 = 1.17e-05  mcm3d_cc_w_0_300_s_1_000 = 5.13e-11  mcm3d_cf_w_0_300_s_1_000 = 5.75e-12
+ mcm3d_ca_w_0_300_s_1_200 = 1.17e-05  mcm3d_cc_w_0_300_s_1_200 = 4.55e-11  mcm3d_cf_w_0_300_s_1_200 = 6.76e-12
+ mcm3d_ca_w_0_300_s_2_100 = 1.17e-05  mcm3d_cc_w_0_300_s_2_100 = 3.06e-11  mcm3d_cf_w_0_300_s_2_100 = 1.12e-11
+ mcm3d_ca_w_0_300_s_3_300 = 1.17e-05  mcm3d_cc_w_0_300_s_3_300 = 2.15e-11  mcm3d_cf_w_0_300_s_3_300 = 1.55e-11
+ mcm3d_ca_w_0_300_s_9_000 = 1.17e-05  mcm3d_cc_w_0_300_s_9_000 = 6.66e-12  mcm3d_cf_w_0_300_s_9_000 = 2.66e-11
+ mcm3d_ca_w_2_400_s_0_300 = 1.17e-05  mcm3d_cc_w_2_400_s_0_300 = 1.17e-10  mcm3d_cf_w_2_400_s_0_300 = 2.02e-12
+ mcm3d_ca_w_2_400_s_0_360 = 1.17e-05  mcm3d_cc_w_2_400_s_0_360 = 1.11e-10  mcm3d_cf_w_2_400_s_0_360 = 2.36e-12
+ mcm3d_ca_w_2_400_s_0_450 = 1.17e-05  mcm3d_cc_w_2_400_s_0_450 = 1.02e-10  mcm3d_cf_w_2_400_s_0_450 = 2.86e-12
+ mcm3d_ca_w_2_400_s_0_600 = 1.17e-05  mcm3d_cc_w_2_400_s_0_600 = 8.93e-11  mcm3d_cf_w_2_400_s_0_600 = 3.69e-12
+ mcm3d_ca_w_2_400_s_0_800 = 1.17e-05  mcm3d_cc_w_2_400_s_0_800 = 7.69e-11  mcm3d_cf_w_2_400_s_0_800 = 4.76e-12
+ mcm3d_ca_w_2_400_s_1_000 = 1.17e-05  mcm3d_cc_w_2_400_s_1_000 = 6.75e-11  mcm3d_cf_w_2_400_s_1_000 = 5.82e-12
+ mcm3d_ca_w_2_400_s_1_200 = 1.17e-05  mcm3d_cc_w_2_400_s_1_200 = 6.04e-11  mcm3d_cf_w_2_400_s_1_200 = 6.85e-12
+ mcm3d_ca_w_2_400_s_2_100 = 1.17e-05  mcm3d_cc_w_2_400_s_2_100 = 4.19e-11  mcm3d_cf_w_2_400_s_2_100 = 1.11e-11
+ mcm3d_ca_w_2_400_s_3_300 = 1.17e-05  mcm3d_cc_w_2_400_s_3_300 = 2.99e-11  mcm3d_cf_w_2_400_s_3_300 = 1.60e-11
+ mcm3d_ca_w_2_400_s_9_000 = 1.17e-05  mcm3d_cc_w_2_400_s_9_000 = 1.04e-11  mcm3d_cf_w_2_400_s_9_000 = 2.94e-11
+ mcm3p1_ca_w_0_300_s_0_300 = 1.26e-05  mcm3p1_cc_w_0_300_s_0_300 = 9.13e-11  mcm3p1_cf_w_0_300_s_0_300 = 2.16e-12
+ mcm3p1_ca_w_0_300_s_0_360 = 1.26e-05  mcm3p1_cc_w_0_300_s_0_360 = 8.60e-11  mcm3p1_cf_w_0_300_s_0_360 = 2.52e-12
+ mcm3p1_ca_w_0_300_s_0_450 = 1.26e-05  mcm3p1_cc_w_0_300_s_0_450 = 7.84e-11  mcm3p1_cf_w_0_300_s_0_450 = 3.09e-12
+ mcm3p1_ca_w_0_300_s_0_600 = 1.26e-05  mcm3p1_cc_w_0_300_s_0_600 = 6.83e-11  mcm3p1_cf_w_0_300_s_0_600 = 4.01e-12
+ mcm3p1_ca_w_0_300_s_0_800 = 1.26e-05  mcm3p1_cc_w_0_300_s_0_800 = 5.83e-11  mcm3p1_cf_w_0_300_s_0_800 = 5.10e-12
+ mcm3p1_ca_w_0_300_s_1_000 = 1.26e-05  mcm3p1_cc_w_0_300_s_1_000 = 5.08e-11  mcm3p1_cf_w_0_300_s_1_000 = 6.21e-12
+ mcm3p1_ca_w_0_300_s_1_200 = 1.26e-05  mcm3p1_cc_w_0_300_s_1_200 = 4.50e-11  mcm3p1_cf_w_0_300_s_1_200 = 7.29e-12
+ mcm3p1_ca_w_0_300_s_2_100 = 1.26e-05  mcm3p1_cc_w_0_300_s_2_100 = 3.00e-11  mcm3p1_cf_w_0_300_s_2_100 = 1.20e-11
+ mcm3p1_ca_w_0_300_s_3_300 = 1.26e-05  mcm3p1_cc_w_0_300_s_3_300 = 2.08e-11  mcm3p1_cf_w_0_300_s_3_300 = 1.65e-11
+ mcm3p1_ca_w_0_300_s_9_000 = 1.26e-05  mcm3p1_cc_w_0_300_s_9_000 = 6.21e-12  mcm3p1_cf_w_0_300_s_9_000 = 2.77e-11
+ mcm3p1_ca_w_2_400_s_0_300 = 1.26e-05  mcm3p1_cc_w_2_400_s_0_300 = 1.16e-10  mcm3p1_cf_w_2_400_s_0_300 = 2.21e-12
+ mcm3p1_ca_w_2_400_s_0_360 = 1.26e-05  mcm3p1_cc_w_2_400_s_0_360 = 1.10e-10  mcm3p1_cf_w_2_400_s_0_360 = 2.58e-12
+ mcm3p1_ca_w_2_400_s_0_450 = 1.26e-05  mcm3p1_cc_w_2_400_s_0_450 = 1.01e-10  mcm3p1_cf_w_2_400_s_0_450 = 3.12e-12
+ mcm3p1_ca_w_2_400_s_0_600 = 1.26e-05  mcm3p1_cc_w_2_400_s_0_600 = 8.83e-11  mcm3p1_cf_w_2_400_s_0_600 = 4.01e-12
+ mcm3p1_ca_w_2_400_s_0_800 = 1.26e-05  mcm3p1_cc_w_2_400_s_0_800 = 7.61e-11  mcm3p1_cf_w_2_400_s_0_800 = 5.17e-12
+ mcm3p1_ca_w_2_400_s_1_000 = 1.26e-05  mcm3p1_cc_w_2_400_s_1_000 = 6.67e-11  mcm3p1_cf_w_2_400_s_1_000 = 6.30e-12
+ mcm3p1_ca_w_2_400_s_1_200 = 1.26e-05  mcm3p1_cc_w_2_400_s_1_200 = 5.96e-11  mcm3p1_cf_w_2_400_s_1_200 = 7.41e-12
+ mcm3p1_ca_w_2_400_s_2_100 = 1.26e-05  mcm3p1_cc_w_2_400_s_2_100 = 4.11e-11  mcm3p1_cf_w_2_400_s_2_100 = 1.20e-11
+ mcm3p1_ca_w_2_400_s_3_300 = 1.26e-05  mcm3p1_cc_w_2_400_s_3_300 = 2.90e-11  mcm3p1_cf_w_2_400_s_3_300 = 1.71e-11
+ mcm3p1_ca_w_2_400_s_9_000 = 1.26e-05  mcm3p1_cc_w_2_400_s_9_000 = 9.88e-12  mcm3p1_cf_w_2_400_s_9_000 = 3.07e-11
+ mcm3l1_ca_w_0_300_s_0_300 = 1.63e-05  mcm3l1_cc_w_0_300_s_0_300 = 9.03e-11  mcm3l1_cf_w_0_300_s_0_300 = 2.77e-12
+ mcm3l1_ca_w_0_300_s_0_360 = 1.63e-05  mcm3l1_cc_w_0_300_s_0_360 = 8.49e-11  mcm3l1_cf_w_0_300_s_0_360 = 3.23e-12
+ mcm3l1_ca_w_0_300_s_0_450 = 1.63e-05  mcm3l1_cc_w_0_300_s_0_450 = 7.73e-11  mcm3l1_cf_w_0_300_s_0_450 = 3.95e-12
+ mcm3l1_ca_w_0_300_s_0_600 = 1.63e-05  mcm3l1_cc_w_0_300_s_0_600 = 6.70e-11  mcm3l1_cf_w_0_300_s_0_600 = 5.10e-12
+ mcm3l1_ca_w_0_300_s_0_800 = 1.63e-05  mcm3l1_cc_w_0_300_s_0_800 = 5.70e-11  mcm3l1_cf_w_0_300_s_0_800 = 6.48e-12
+ mcm3l1_ca_w_0_300_s_1_000 = 1.63e-05  mcm3l1_cc_w_0_300_s_1_000 = 4.93e-11  mcm3l1_cf_w_0_300_s_1_000 = 7.87e-12
+ mcm3l1_ca_w_0_300_s_1_200 = 1.63e-05  mcm3l1_cc_w_0_300_s_1_200 = 4.33e-11  mcm3l1_cf_w_0_300_s_1_200 = 9.21e-12
+ mcm3l1_ca_w_0_300_s_2_100 = 1.63e-05  mcm3l1_cc_w_0_300_s_2_100 = 2.79e-11  mcm3l1_cf_w_0_300_s_2_100 = 1.49e-11
+ mcm3l1_ca_w_0_300_s_3_300 = 1.63e-05  mcm3l1_cc_w_0_300_s_3_300 = 1.87e-11  mcm3l1_cf_w_0_300_s_3_300 = 2.00e-11
+ mcm3l1_ca_w_0_300_s_9_000 = 1.63e-05  mcm3l1_cc_w_0_300_s_9_000 = 5.07e-12  mcm3l1_cf_w_0_300_s_9_000 = 3.11e-11
+ mcm3l1_ca_w_2_400_s_0_300 = 1.63e-05  mcm3l1_cc_w_2_400_s_0_300 = 1.14e-10  mcm3l1_cf_w_2_400_s_0_300 = 2.80e-12
+ mcm3l1_ca_w_2_400_s_0_360 = 1.63e-05  mcm3l1_cc_w_2_400_s_0_360 = 1.07e-10  mcm3l1_cf_w_2_400_s_0_360 = 3.26e-12
+ mcm3l1_ca_w_2_400_s_0_450 = 1.63e-05  mcm3l1_cc_w_2_400_s_0_450 = 9.83e-11  mcm3l1_cf_w_2_400_s_0_450 = 3.95e-12
+ mcm3l1_ca_w_2_400_s_0_600 = 1.63e-05  mcm3l1_cc_w_2_400_s_0_600 = 8.58e-11  mcm3l1_cf_w_2_400_s_0_600 = 5.08e-12
+ mcm3l1_ca_w_2_400_s_0_800 = 1.63e-05  mcm3l1_cc_w_2_400_s_0_800 = 7.35e-11  mcm3l1_cf_w_2_400_s_0_800 = 6.54e-12
+ mcm3l1_ca_w_2_400_s_1_000 = 1.63e-05  mcm3l1_cc_w_2_400_s_1_000 = 6.40e-11  mcm3l1_cf_w_2_400_s_1_000 = 7.95e-12
+ mcm3l1_ca_w_2_400_s_1_200 = 1.63e-05  mcm3l1_cc_w_2_400_s_1_200 = 5.69e-11  mcm3l1_cf_w_2_400_s_1_200 = 9.31e-12
+ mcm3l1_ca_w_2_400_s_2_100 = 1.63e-05  mcm3l1_cc_w_2_400_s_2_100 = 3.84e-11  mcm3l1_cf_w_2_400_s_2_100 = 1.48e-11
+ mcm3l1_ca_w_2_400_s_3_300 = 1.63e-05  mcm3l1_cc_w_2_400_s_3_300 = 2.66e-11  mcm3l1_cf_w_2_400_s_3_300 = 2.08e-11
+ mcm3l1_ca_w_2_400_s_9_000 = 1.63e-05  mcm3l1_cc_w_2_400_s_9_000 = 8.40e-12  mcm3l1_cf_w_2_400_s_9_000 = 3.46e-11
+ mcm3m1_ca_w_0_300_s_0_300 = 2.58e-05  mcm3m1_cc_w_0_300_s_0_300 = 8.82e-11  mcm3m1_cf_w_0_300_s_0_300 = 4.30e-12
+ mcm3m1_ca_w_0_300_s_0_360 = 2.58e-05  mcm3m1_cc_w_0_300_s_0_360 = 8.25e-11  mcm3m1_cf_w_0_300_s_0_360 = 5.01e-12
+ mcm3m1_ca_w_0_300_s_0_450 = 2.58e-05  mcm3m1_cc_w_0_300_s_0_450 = 7.47e-11  mcm3m1_cf_w_0_300_s_0_450 = 6.08e-12
+ mcm3m1_ca_w_0_300_s_0_600 = 2.58e-05  mcm3m1_cc_w_0_300_s_0_600 = 6.42e-11  mcm3m1_cf_w_0_300_s_0_600 = 7.80e-12
+ mcm3m1_ca_w_0_300_s_0_800 = 2.58e-05  mcm3m1_cc_w_0_300_s_0_800 = 5.39e-11  mcm3m1_cf_w_0_300_s_0_800 = 9.84e-12
+ mcm3m1_ca_w_0_300_s_1_000 = 2.58e-05  mcm3m1_cc_w_0_300_s_1_000 = 4.59e-11  mcm3m1_cf_w_0_300_s_1_000 = 1.18e-11
+ mcm3m1_ca_w_0_300_s_1_200 = 2.58e-05  mcm3m1_cc_w_0_300_s_1_200 = 3.99e-11  mcm3m1_cf_w_0_300_s_1_200 = 1.37e-11
+ mcm3m1_ca_w_0_300_s_2_100 = 2.58e-05  mcm3m1_cc_w_0_300_s_2_100 = 2.40e-11  mcm3m1_cf_w_0_300_s_2_100 = 2.13e-11
+ mcm3m1_ca_w_0_300_s_3_300 = 2.58e-05  mcm3m1_cc_w_0_300_s_3_300 = 1.51e-11  mcm3m1_cf_w_0_300_s_3_300 = 2.72e-11
+ mcm3m1_ca_w_0_300_s_9_000 = 2.58e-05  mcm3m1_cc_w_0_300_s_9_000 = 3.46e-12  mcm3m1_cf_w_0_300_s_9_000 = 3.75e-11
+ mcm3m1_ca_w_2_400_s_0_300 = 2.58e-05  mcm3m1_cc_w_2_400_s_0_300 = 1.09e-10  mcm3m1_cf_w_2_400_s_0_300 = 4.32e-12
+ mcm3m1_ca_w_2_400_s_0_360 = 2.58e-05  mcm3m1_cc_w_2_400_s_0_360 = 1.02e-10  mcm3m1_cf_w_2_400_s_0_360 = 5.03e-12
+ mcm3m1_ca_w_2_400_s_0_450 = 2.58e-05  mcm3m1_cc_w_2_400_s_0_450 = 9.35e-11  mcm3m1_cf_w_2_400_s_0_450 = 6.07e-12
+ mcm3m1_ca_w_2_400_s_0_600 = 2.58e-05  mcm3m1_cc_w_2_400_s_0_600 = 8.09e-11  mcm3m1_cf_w_2_400_s_0_600 = 7.76e-12
+ mcm3m1_ca_w_2_400_s_0_800 = 2.58e-05  mcm3m1_cc_w_2_400_s_0_800 = 6.86e-11  mcm3m1_cf_w_2_400_s_0_800 = 9.91e-12
+ mcm3m1_ca_w_2_400_s_1_000 = 2.58e-05  mcm3m1_cc_w_2_400_s_1_000 = 5.93e-11  mcm3m1_cf_w_2_400_s_1_000 = 1.20e-11
+ mcm3m1_ca_w_2_400_s_1_200 = 2.58e-05  mcm3m1_cc_w_2_400_s_1_200 = 5.22e-11  mcm3m1_cf_w_2_400_s_1_200 = 1.39e-11
+ mcm3m1_ca_w_2_400_s_2_100 = 2.58e-05  mcm3m1_cc_w_2_400_s_2_100 = 3.39e-11  mcm3m1_cf_w_2_400_s_2_100 = 2.12e-11
+ mcm3m1_ca_w_2_400_s_3_300 = 2.58e-05  mcm3m1_cc_w_2_400_s_3_300 = 2.24e-11  mcm3m1_cf_w_2_400_s_3_300 = 2.83e-11
+ mcm3m1_ca_w_2_400_s_9_000 = 2.58e-05  mcm3m1_cc_w_2_400_s_9_000 = 6.40e-12  mcm3m1_cf_w_2_400_s_9_000 = 4.19e-11
+ mcm3m2_ca_w_0_300_s_0_300 = 5.95e-05  mcm3m2_cc_w_0_300_s_0_300 = 8.18e-11  mcm3m2_cf_w_0_300_s_0_300 = 9.43e-12
+ mcm3m2_ca_w_0_300_s_0_360 = 5.95e-05  mcm3m2_cc_w_0_300_s_0_360 = 7.61e-11  mcm3m2_cf_w_0_300_s_0_360 = 1.09e-11
+ mcm3m2_ca_w_0_300_s_0_450 = 5.95e-05  mcm3m2_cc_w_0_300_s_0_450 = 6.80e-11  mcm3m2_cf_w_0_300_s_0_450 = 1.30e-11
+ mcm3m2_ca_w_0_300_s_0_600 = 5.95e-05  mcm3m2_cc_w_0_300_s_0_600 = 5.72e-11  mcm3m2_cf_w_0_300_s_0_600 = 1.63e-11
+ mcm3m2_ca_w_0_300_s_0_800 = 5.95e-05  mcm3m2_cc_w_0_300_s_0_800 = 4.66e-11  mcm3m2_cf_w_0_300_s_0_800 = 2.00e-11
+ mcm3m2_ca_w_0_300_s_1_000 = 5.95e-05  mcm3m2_cc_w_0_300_s_1_000 = 3.86e-11  mcm3m2_cf_w_0_300_s_1_000 = 2.34e-11
+ mcm3m2_ca_w_0_300_s_1_200 = 5.95e-05  mcm3m2_cc_w_0_300_s_1_200 = 3.25e-11  mcm3m2_cf_w_0_300_s_1_200 = 2.63e-11
+ mcm3m2_ca_w_0_300_s_2_100 = 5.95e-05  mcm3m2_cc_w_0_300_s_2_100 = 1.73e-11  mcm3m2_cf_w_0_300_s_2_100 = 3.64e-11
+ mcm3m2_ca_w_0_300_s_3_300 = 5.95e-05  mcm3m2_cc_w_0_300_s_3_300 = 9.90e-12  mcm3m2_cf_w_0_300_s_3_300 = 4.26e-11
+ mcm3m2_ca_w_0_300_s_9_000 = 5.95e-05  mcm3m2_cc_w_0_300_s_9_000 = 2.00e-12  mcm3m2_cf_w_0_300_s_9_000 = 5.01e-11
+ mcm3m2_ca_w_2_400_s_0_300 = 5.95e-05  mcm3m2_cc_w_2_400_s_0_300 = 9.95e-11  mcm3m2_cf_w_2_400_s_0_300 = 9.45e-12
+ mcm3m2_ca_w_2_400_s_0_360 = 5.95e-05  mcm3m2_cc_w_2_400_s_0_360 = 9.32e-11  mcm3m2_cf_w_2_400_s_0_360 = 1.09e-11
+ mcm3m2_ca_w_2_400_s_0_450 = 5.95e-05  mcm3m2_cc_w_2_400_s_0_450 = 8.42e-11  mcm3m2_cf_w_2_400_s_0_450 = 1.30e-11
+ mcm3m2_ca_w_2_400_s_0_600 = 5.95e-05  mcm3m2_cc_w_2_400_s_0_600 = 7.22e-11  mcm3m2_cf_w_2_400_s_0_600 = 1.62e-11
+ mcm3m2_ca_w_2_400_s_0_800 = 5.95e-05  mcm3m2_cc_w_2_400_s_0_800 = 6.00e-11  mcm3m2_cf_w_2_400_s_0_800 = 2.01e-11
+ mcm3m2_ca_w_2_400_s_1_000 = 5.95e-05  mcm3m2_cc_w_2_400_s_1_000 = 5.08e-11  mcm3m2_cf_w_2_400_s_1_000 = 2.35e-11
+ mcm3m2_ca_w_2_400_s_1_200 = 5.95e-05  mcm3m2_cc_w_2_400_s_1_200 = 4.41e-11  mcm3m2_cf_w_2_400_s_1_200 = 2.65e-11
+ mcm3m2_ca_w_2_400_s_2_100 = 5.95e-05  mcm3m2_cc_w_2_400_s_2_100 = 2.70e-11  mcm3m2_cf_w_2_400_s_2_100 = 3.65e-11
+ mcm3m2_ca_w_2_400_s_3_300 = 5.95e-05  mcm3m2_cc_w_2_400_s_3_300 = 1.69e-11  mcm3m2_cf_w_2_400_s_3_300 = 4.44e-11
+ mcm3m2_ca_w_2_400_s_9_000 = 5.95e-05  mcm3m2_cc_w_2_400_s_9_000 = 4.35e-12  mcm3m2_cf_w_2_400_s_9_000 = 5.60e-11
+ mcm4f_ca_w_0_300_s_0_300 = 7.28e-06  mcm4f_cc_w_0_300_s_0_300 = 9.29e-11  mcm4f_cf_w_0_300_s_0_300 = 1.25e-12
+ mcm4f_ca_w_0_300_s_0_360 = 7.28e-06  mcm4f_cc_w_0_300_s_0_360 = 8.74e-11  mcm4f_cf_w_0_300_s_0_360 = 1.46e-12
+ mcm4f_ca_w_0_300_s_0_450 = 7.28e-06  mcm4f_cc_w_0_300_s_0_450 = 8.02e-11  mcm4f_cf_w_0_300_s_0_450 = 1.80e-12
+ mcm4f_ca_w_0_300_s_0_600 = 7.28e-06  mcm4f_cc_w_0_300_s_0_600 = 7.04e-11  mcm4f_cf_w_0_300_s_0_600 = 2.36e-12
+ mcm4f_ca_w_0_300_s_0_800 = 7.28e-06  mcm4f_cc_w_0_300_s_0_800 = 6.10e-11  mcm4f_cf_w_0_300_s_0_800 = 3.00e-12
+ mcm4f_ca_w_0_300_s_1_000 = 7.28e-06  mcm4f_cc_w_0_300_s_1_000 = 5.37e-11  mcm4f_cf_w_0_300_s_1_000 = 3.66e-12
+ mcm4f_ca_w_0_300_s_1_200 = 7.28e-06  mcm4f_cc_w_0_300_s_1_200 = 4.82e-11  mcm4f_cf_w_0_300_s_1_200 = 4.32e-12
+ mcm4f_ca_w_0_300_s_2_100 = 7.28e-06  mcm4f_cc_w_0_300_s_2_100 = 3.39e-11  mcm4f_cf_w_0_300_s_2_100 = 7.40e-12
+ mcm4f_ca_w_0_300_s_3_300 = 7.28e-06  mcm4f_cc_w_0_300_s_3_300 = 2.51e-11  mcm4f_cf_w_0_300_s_3_300 = 1.05e-11
+ mcm4f_ca_w_0_300_s_9_000 = 7.28e-06  mcm4f_cc_w_0_300_s_9_000 = 9.35e-12  mcm4f_cf_w_0_300_s_9_000 = 2.04e-11
+ mcm4f_ca_w_2_400_s_0_300 = 7.28e-06  mcm4f_cc_w_2_400_s_0_300 = 1.21e-10  mcm4f_cf_w_2_400_s_0_300 = 1.26e-12
+ mcm4f_ca_w_2_400_s_0_360 = 7.28e-06  mcm4f_cc_w_2_400_s_0_360 = 1.15e-10  mcm4f_cf_w_2_400_s_0_360 = 1.48e-12
+ mcm4f_ca_w_2_400_s_0_450 = 7.28e-06  mcm4f_cc_w_2_400_s_0_450 = 1.06e-10  mcm4f_cf_w_2_400_s_0_450 = 1.80e-12
+ mcm4f_ca_w_2_400_s_0_600 = 7.28e-06  mcm4f_cc_w_2_400_s_0_600 = 9.38e-11  mcm4f_cf_w_2_400_s_0_600 = 2.32e-12
+ mcm4f_ca_w_2_400_s_0_800 = 7.28e-06  mcm4f_cc_w_2_400_s_0_800 = 8.14e-11  mcm4f_cf_w_2_400_s_0_800 = 3.02e-12
+ mcm4f_ca_w_2_400_s_1_000 = 7.28e-06  mcm4f_cc_w_2_400_s_1_000 = 7.20e-11  mcm4f_cf_w_2_400_s_1_000 = 3.71e-12
+ mcm4f_ca_w_2_400_s_1_200 = 7.28e-06  mcm4f_cc_w_2_400_s_1_200 = 6.49e-11  mcm4f_cf_w_2_400_s_1_200 = 4.37e-12
+ mcm4f_ca_w_2_400_s_2_100 = 7.28e-06  mcm4f_cc_w_2_400_s_2_100 = 4.64e-11  mcm4f_cf_w_2_400_s_2_100 = 7.27e-12
+ mcm4f_ca_w_2_400_s_3_300 = 7.28e-06  mcm4f_cc_w_2_400_s_3_300 = 3.42e-11  mcm4f_cf_w_2_400_s_3_300 = 1.08e-11
+ mcm4f_ca_w_2_400_s_9_000 = 7.28e-06  mcm4f_cc_w_2_400_s_9_000 = 1.36e-11  mcm4f_cf_w_2_400_s_9_000 = 2.23e-11
+ mcm4d_ca_w_0_300_s_0_300 = 7.98e-06  mcm4d_cc_w_0_300_s_0_300 = 9.27e-11  mcm4d_cf_w_0_300_s_0_300 = 1.37e-12
+ mcm4d_ca_w_0_300_s_0_360 = 7.98e-06  mcm4d_cc_w_0_300_s_0_360 = 8.72e-11  mcm4d_cf_w_0_300_s_0_360 = 1.60e-12
+ mcm4d_ca_w_0_300_s_0_450 = 7.98e-06  mcm4d_cc_w_0_300_s_0_450 = 8.00e-11  mcm4d_cf_w_0_300_s_0_450 = 1.97e-12
+ mcm4d_ca_w_0_300_s_0_600 = 7.98e-06  mcm4d_cc_w_0_300_s_0_600 = 7.02e-11  mcm4d_cf_w_0_300_s_0_600 = 2.57e-12
+ mcm4d_ca_w_0_300_s_0_800 = 7.98e-06  mcm4d_cc_w_0_300_s_0_800 = 6.08e-11  mcm4d_cf_w_0_300_s_0_800 = 3.27e-12
+ mcm4d_ca_w_0_300_s_1_000 = 7.98e-06  mcm4d_cc_w_0_300_s_1_000 = 5.34e-11  mcm4d_cf_w_0_300_s_1_000 = 3.99e-12
+ mcm4d_ca_w_0_300_s_1_200 = 7.98e-06  mcm4d_cc_w_0_300_s_1_200 = 4.78e-11  mcm4d_cf_w_0_300_s_1_200 = 4.72e-12
+ mcm4d_ca_w_0_300_s_2_100 = 7.98e-06  mcm4d_cc_w_0_300_s_2_100 = 3.33e-11  mcm4d_cf_w_0_300_s_2_100 = 8.03e-12
+ mcm4d_ca_w_0_300_s_3_300 = 7.98e-06  mcm4d_cc_w_0_300_s_3_300 = 2.44e-11  mcm4d_cf_w_0_300_s_3_300 = 1.13e-11
+ mcm4d_ca_w_0_300_s_9_000 = 7.98e-06  mcm4d_cc_w_0_300_s_9_000 = 8.75e-12  mcm4d_cf_w_0_300_s_9_000 = 2.16e-11
+ mcm4d_ca_w_2_400_s_0_300 = 7.98e-06  mcm4d_cc_w_2_400_s_0_300 = 1.21e-10  mcm4d_cf_w_2_400_s_0_300 = 1.39e-12
+ mcm4d_ca_w_2_400_s_0_360 = 7.98e-06  mcm4d_cc_w_2_400_s_0_360 = 1.14e-10  mcm4d_cf_w_2_400_s_0_360 = 1.62e-12
+ mcm4d_ca_w_2_400_s_0_450 = 7.98e-06  mcm4d_cc_w_2_400_s_0_450 = 1.05e-10  mcm4d_cf_w_2_400_s_0_450 = 1.97e-12
+ mcm4d_ca_w_2_400_s_0_600 = 7.98e-06  mcm4d_cc_w_2_400_s_0_600 = 9.31e-11  mcm4d_cf_w_2_400_s_0_600 = 2.55e-12
+ mcm4d_ca_w_2_400_s_0_800 = 7.98e-06  mcm4d_cc_w_2_400_s_0_800 = 8.07e-11  mcm4d_cf_w_2_400_s_0_800 = 3.30e-12
+ mcm4d_ca_w_2_400_s_1_000 = 7.98e-06  mcm4d_cc_w_2_400_s_1_000 = 7.13e-11  mcm4d_cf_w_2_400_s_1_000 = 4.04e-12
+ mcm4d_ca_w_2_400_s_1_200 = 7.98e-06  mcm4d_cc_w_2_400_s_1_200 = 6.41e-11  mcm4d_cf_w_2_400_s_1_200 = 4.77e-12
+ mcm4d_ca_w_2_400_s_2_100 = 7.98e-06  mcm4d_cc_w_2_400_s_2_100 = 4.55e-11  mcm4d_cf_w_2_400_s_2_100 = 7.90e-12
+ mcm4d_ca_w_2_400_s_3_300 = 7.98e-06  mcm4d_cc_w_2_400_s_3_300 = 3.33e-11  mcm4d_cf_w_2_400_s_3_300 = 1.16e-11
+ mcm4d_ca_w_2_400_s_9_000 = 7.98e-06  mcm4d_cc_w_2_400_s_9_000 = 1.29e-11  mcm4d_cf_w_2_400_s_9_000 = 2.36e-11
+ mcm4p1_ca_w_0_300_s_0_300 = 8.42e-06  mcm4p1_cc_w_0_300_s_0_300 = 9.26e-11  mcm4p1_cf_w_0_300_s_0_300 = 1.45e-12
+ mcm4p1_ca_w_0_300_s_0_360 = 8.42e-06  mcm4p1_cc_w_0_300_s_0_360 = 8.72e-11  mcm4p1_cf_w_0_300_s_0_360 = 1.69e-12
+ mcm4p1_ca_w_0_300_s_0_450 = 8.42e-06  mcm4p1_cc_w_0_300_s_0_450 = 7.99e-11  mcm4p1_cf_w_0_300_s_0_450 = 2.08e-12
+ mcm4p1_ca_w_0_300_s_0_600 = 8.42e-06  mcm4p1_cc_w_0_300_s_0_600 = 7.00e-11  mcm4p1_cf_w_0_300_s_0_600 = 2.72e-12
+ mcm4p1_ca_w_0_300_s_0_800 = 8.42e-06  mcm4p1_cc_w_0_300_s_0_800 = 6.05e-11  mcm4p1_cf_w_0_300_s_0_800 = 3.45e-12
+ mcm4p1_ca_w_0_300_s_1_000 = 8.42e-06  mcm4p1_cc_w_0_300_s_1_000 = 5.31e-11  mcm4p1_cf_w_0_300_s_1_000 = 4.21e-12
+ mcm4p1_ca_w_0_300_s_1_200 = 8.42e-06  mcm4p1_cc_w_0_300_s_1_200 = 4.75e-11  mcm4p1_cf_w_0_300_s_1_200 = 4.97e-12
+ mcm4p1_ca_w_0_300_s_2_100 = 8.42e-06  mcm4p1_cc_w_0_300_s_2_100 = 3.30e-11  mcm4p1_cf_w_0_300_s_2_100 = 8.42e-12
+ mcm4p1_ca_w_0_300_s_3_300 = 8.42e-06  mcm4p1_cc_w_0_300_s_3_300 = 2.40e-11  mcm4p1_cf_w_0_300_s_3_300 = 1.18e-11
+ mcm4p1_ca_w_0_300_s_9_000 = 8.42e-06  mcm4p1_cc_w_0_300_s_9_000 = 8.39e-12  mcm4p1_cf_w_0_300_s_9_000 = 2.23e-11
+ mcm4p1_ca_w_2_400_s_0_300 = 8.42e-06  mcm4p1_cc_w_2_400_s_0_300 = 1.20e-10  mcm4p1_cf_w_2_400_s_0_300 = 1.48e-12
+ mcm4p1_ca_w_2_400_s_0_360 = 8.42e-06  mcm4p1_cc_w_2_400_s_0_360 = 1.14e-10  mcm4p1_cf_w_2_400_s_0_360 = 1.72e-12
+ mcm4p1_ca_w_2_400_s_0_450 = 8.42e-06  mcm4p1_cc_w_2_400_s_0_450 = 1.05e-10  mcm4p1_cf_w_2_400_s_0_450 = 2.09e-12
+ mcm4p1_ca_w_2_400_s_0_600 = 8.42e-06  mcm4p1_cc_w_2_400_s_0_600 = 9.25e-11  mcm4p1_cf_w_2_400_s_0_600 = 2.70e-12
+ mcm4p1_ca_w_2_400_s_0_800 = 8.42e-06  mcm4p1_cc_w_2_400_s_0_800 = 8.03e-11  mcm4p1_cf_w_2_400_s_0_800 = 3.49e-12
+ mcm4p1_ca_w_2_400_s_1_000 = 8.42e-06  mcm4p1_cc_w_2_400_s_1_000 = 7.08e-11  mcm4p1_cf_w_2_400_s_1_000 = 4.27e-12
+ mcm4p1_ca_w_2_400_s_1_200 = 8.42e-06  mcm4p1_cc_w_2_400_s_1_200 = 6.37e-11  mcm4p1_cf_w_2_400_s_1_200 = 5.04e-12
+ mcm4p1_ca_w_2_400_s_2_100 = 8.42e-06  mcm4p1_cc_w_2_400_s_2_100 = 4.50e-11  mcm4p1_cf_w_2_400_s_2_100 = 8.31e-12
+ mcm4p1_ca_w_2_400_s_3_300 = 8.42e-06  mcm4p1_cc_w_2_400_s_3_300 = 3.28e-11  mcm4p1_cf_w_2_400_s_3_300 = 1.22e-11
+ mcm4p1_ca_w_2_400_s_9_000 = 8.42e-06  mcm4p1_cc_w_2_400_s_9_000 = 1.24e-11  mcm4p1_cf_w_2_400_s_9_000 = 2.45e-11
+ mcm4l1_ca_w_0_300_s_0_300 = 9.92e-06  mcm4l1_cc_w_0_300_s_0_300 = 9.22e-11  mcm4l1_cf_w_0_300_s_0_300 = 1.70e-12
+ mcm4l1_ca_w_0_300_s_0_360 = 9.92e-06  mcm4l1_cc_w_0_300_s_0_360 = 8.68e-11  mcm4l1_cf_w_0_300_s_0_360 = 1.99e-12
+ mcm4l1_ca_w_0_300_s_0_450 = 9.92e-06  mcm4l1_cc_w_0_300_s_0_450 = 7.94e-11  mcm4l1_cf_w_0_300_s_0_450 = 2.44e-12
+ mcm4l1_ca_w_0_300_s_0_600 = 9.92e-06  mcm4l1_cc_w_0_300_s_0_600 = 6.95e-11  mcm4l1_cf_w_0_300_s_0_600 = 3.18e-12
+ mcm4l1_ca_w_0_300_s_0_800 = 9.92e-06  mcm4l1_cc_w_0_300_s_0_800 = 5.99e-11  mcm4l1_cf_w_0_300_s_0_800 = 4.03e-12
+ mcm4l1_ca_w_0_300_s_1_000 = 9.92e-06  mcm4l1_cc_w_0_300_s_1_000 = 5.24e-11  mcm4l1_cf_w_0_300_s_1_000 = 4.91e-12
+ mcm4l1_ca_w_0_300_s_1_200 = 9.92e-06  mcm4l1_cc_w_0_300_s_1_200 = 4.67e-11  mcm4l1_cf_w_0_300_s_1_200 = 5.80e-12
+ mcm4l1_ca_w_0_300_s_2_100 = 9.92e-06  mcm4l1_cc_w_0_300_s_2_100 = 3.20e-11  mcm4l1_cf_w_0_300_s_2_100 = 9.72e-12
+ mcm4l1_ca_w_0_300_s_3_300 = 9.92e-06  mcm4l1_cc_w_0_300_s_3_300 = 2.28e-11  mcm4l1_cf_w_0_300_s_3_300 = 1.36e-11
+ mcm4l1_ca_w_0_300_s_9_000 = 9.92e-06  mcm4l1_cc_w_0_300_s_9_000 = 7.41e-12  mcm4l1_cf_w_0_300_s_9_000 = 2.44e-11
+ mcm4l1_ca_w_2_400_s_0_300 = 9.92e-06  mcm4l1_cc_w_2_400_s_0_300 = 1.19e-10  mcm4l1_cf_w_2_400_s_0_300 = 1.71e-12
+ mcm4l1_ca_w_2_400_s_0_360 = 9.92e-06  mcm4l1_cc_w_2_400_s_0_360 = 1.13e-10  mcm4l1_cf_w_2_400_s_0_360 = 2.00e-12
+ mcm4l1_ca_w_2_400_s_0_450 = 9.92e-06  mcm4l1_cc_w_2_400_s_0_450 = 1.03e-10  mcm4l1_cf_w_2_400_s_0_450 = 2.43e-12
+ mcm4l1_ca_w_2_400_s_0_600 = 9.92e-06  mcm4l1_cc_w_2_400_s_0_600 = 9.12e-11  mcm4l1_cf_w_2_400_s_0_600 = 3.14e-12
+ mcm4l1_ca_w_2_400_s_0_800 = 9.92e-06  mcm4l1_cc_w_2_400_s_0_800 = 7.88e-11  mcm4l1_cf_w_2_400_s_0_800 = 4.07e-12
+ mcm4l1_ca_w_2_400_s_1_000 = 9.92e-06  mcm4l1_cc_w_2_400_s_1_000 = 6.94e-11  mcm4l1_cf_w_2_400_s_1_000 = 4.97e-12
+ mcm4l1_ca_w_2_400_s_1_200 = 9.92e-06  mcm4l1_cc_w_2_400_s_1_200 = 6.22e-11  mcm4l1_cf_w_2_400_s_1_200 = 5.86e-12
+ mcm4l1_ca_w_2_400_s_2_100 = 9.92e-06  mcm4l1_cc_w_2_400_s_2_100 = 4.35e-11  mcm4l1_cf_w_2_400_s_2_100 = 9.62e-12
+ mcm4l1_ca_w_2_400_s_3_300 = 9.92e-06  mcm4l1_cc_w_2_400_s_3_300 = 3.12e-11  mcm4l1_cf_w_2_400_s_3_300 = 1.40e-11
+ mcm4l1_ca_w_2_400_s_9_000 = 9.92e-06  mcm4l1_cc_w_2_400_s_9_000 = 1.12e-11  mcm4l1_cf_w_2_400_s_9_000 = 2.69e-11
+ mcm4m1_ca_w_0_300_s_0_300 = 1.28e-05  mcm4m1_cc_w_0_300_s_0_300 = 9.15e-11  mcm4m1_cf_w_0_300_s_0_300 = 2.17e-12
+ mcm4m1_ca_w_0_300_s_0_360 = 1.28e-05  mcm4m1_cc_w_0_300_s_0_360 = 8.61e-11  mcm4m1_cf_w_0_300_s_0_360 = 2.54e-12
+ mcm4m1_ca_w_0_300_s_0_450 = 1.28e-05  mcm4m1_cc_w_0_300_s_0_450 = 7.86e-11  mcm4m1_cf_w_0_300_s_0_450 = 3.11e-12
+ mcm4m1_ca_w_0_300_s_0_600 = 1.28e-05  mcm4m1_cc_w_0_300_s_0_600 = 6.85e-11  mcm4m1_cf_w_0_300_s_0_600 = 4.04e-12
+ mcm4m1_ca_w_0_300_s_0_800 = 1.28e-05  mcm4m1_cc_w_0_300_s_0_800 = 5.88e-11  mcm4m1_cf_w_0_300_s_0_800 = 5.13e-12
+ mcm4m1_ca_w_0_300_s_1_000 = 1.28e-05  mcm4m1_cc_w_0_300_s_1_000 = 5.12e-11  mcm4m1_cf_w_0_300_s_1_000 = 6.24e-12
+ mcm4m1_ca_w_0_300_s_1_200 = 1.28e-05  mcm4m1_cc_w_0_300_s_1_200 = 4.54e-11  mcm4m1_cf_w_0_300_s_1_200 = 7.33e-12
+ mcm4m1_ca_w_0_300_s_2_100 = 1.28e-05  mcm4m1_cc_w_0_300_s_2_100 = 3.01e-11  mcm4m1_cf_w_0_300_s_2_100 = 1.21e-11
+ mcm4m1_ca_w_0_300_s_3_300 = 1.28e-05  mcm4m1_cc_w_0_300_s_3_300 = 2.08e-11  mcm4m1_cf_w_0_300_s_3_300 = 1.66e-11
+ mcm4m1_ca_w_0_300_s_9_000 = 1.28e-05  mcm4m1_cc_w_0_300_s_9_000 = 6.00e-12  mcm4m1_cf_w_0_300_s_9_000 = 2.78e-11
+ mcm4m1_ca_w_2_400_s_0_300 = 1.28e-05  mcm4m1_cc_w_2_400_s_0_300 = 1.17e-10  mcm4m1_cf_w_2_400_s_0_300 = 2.18e-12
+ mcm4m1_ca_w_2_400_s_0_360 = 1.28e-05  mcm4m1_cc_w_2_400_s_0_360 = 1.10e-10  mcm4m1_cf_w_2_400_s_0_360 = 2.55e-12
+ mcm4m1_ca_w_2_400_s_0_450 = 1.28e-05  mcm4m1_cc_w_2_400_s_0_450 = 1.01e-10  mcm4m1_cf_w_2_400_s_0_450 = 3.09e-12
+ mcm4m1_ca_w_2_400_s_0_600 = 1.28e-05  mcm4m1_cc_w_2_400_s_0_600 = 8.88e-11  mcm4m1_cf_w_2_400_s_0_600 = 3.99e-12
+ mcm4m1_ca_w_2_400_s_0_800 = 1.28e-05  mcm4m1_cc_w_2_400_s_0_800 = 7.64e-11  mcm4m1_cf_w_2_400_s_0_800 = 5.16e-12
+ mcm4m1_ca_w_2_400_s_1_000 = 1.28e-05  mcm4m1_cc_w_2_400_s_1_000 = 6.70e-11  mcm4m1_cf_w_2_400_s_1_000 = 6.30e-12
+ mcm4m1_ca_w_2_400_s_1_200 = 1.28e-05  mcm4m1_cc_w_2_400_s_1_200 = 5.97e-11  mcm4m1_cf_w_2_400_s_1_200 = 7.40e-12
+ mcm4m1_ca_w_2_400_s_2_100 = 1.28e-05  mcm4m1_cc_w_2_400_s_2_100 = 4.09e-11  mcm4m1_cf_w_2_400_s_2_100 = 1.20e-11
+ mcm4m1_ca_w_2_400_s_3_300 = 1.28e-05  mcm4m1_cc_w_2_400_s_3_300 = 2.87e-11  mcm4m1_cf_w_2_400_s_3_300 = 1.72e-11
+ mcm4m1_ca_w_2_400_s_9_000 = 1.28e-05  mcm4m1_cc_w_2_400_s_9_000 = 9.48e-12  mcm4m1_cf_w_2_400_s_9_000 = 3.08e-11
+ mcm4m2_ca_w_0_300_s_0_300 = 1.78e-05  mcm4m2_cc_w_0_300_s_0_300 = 9.02e-11  mcm4m2_cf_w_0_300_s_0_300 = 3.00e-12
+ mcm4m2_ca_w_0_300_s_0_360 = 1.78e-05  mcm4m2_cc_w_0_300_s_0_360 = 8.48e-11  mcm4m2_cf_w_0_300_s_0_360 = 3.50e-12
+ mcm4m2_ca_w_0_300_s_0_450 = 1.78e-05  mcm4m2_cc_w_0_300_s_0_450 = 7.71e-11  mcm4m2_cf_w_0_300_s_0_450 = 4.27e-12
+ mcm4m2_ca_w_0_300_s_0_600 = 1.78e-05  mcm4m2_cc_w_0_300_s_0_600 = 6.68e-11  mcm4m2_cf_w_0_300_s_0_600 = 5.52e-12
+ mcm4m2_ca_w_0_300_s_0_800 = 1.78e-05  mcm4m2_cc_w_0_300_s_0_800 = 5.69e-11  mcm4m2_cf_w_0_300_s_0_800 = 6.99e-12
+ mcm4m2_ca_w_0_300_s_1_000 = 1.78e-05  mcm4m2_cc_w_0_300_s_1_000 = 4.90e-11  mcm4m2_cf_w_0_300_s_1_000 = 8.47e-12
+ mcm4m2_ca_w_0_300_s_1_200 = 1.78e-05  mcm4m2_cc_w_0_300_s_1_200 = 4.31e-11  mcm4m2_cf_w_0_300_s_1_200 = 9.89e-12
+ mcm4m2_ca_w_0_300_s_2_100 = 1.78e-05  mcm4m2_cc_w_0_300_s_2_100 = 2.75e-11  mcm4m2_cf_w_0_300_s_2_100 = 1.59e-11
+ mcm4m2_ca_w_0_300_s_3_300 = 1.78e-05  mcm4m2_cc_w_0_300_s_3_300 = 1.81e-11  mcm4m2_cf_w_0_300_s_3_300 = 2.12e-11
+ mcm4m2_ca_w_0_300_s_9_000 = 1.78e-05  mcm4m2_cc_w_0_300_s_9_000 = 4.58e-12  mcm4m2_cf_w_0_300_s_9_000 = 3.23e-11
+ mcm4m2_ca_w_2_400_s_0_300 = 1.78e-05  mcm4m2_cc_w_2_400_s_0_300 = 1.13e-10  mcm4m2_cf_w_2_400_s_0_300 = 3.01e-12
+ mcm4m2_ca_w_2_400_s_0_360 = 1.78e-05  mcm4m2_cc_w_2_400_s_0_360 = 1.07e-10  mcm4m2_cf_w_2_400_s_0_360 = 3.51e-12
+ mcm4m2_ca_w_2_400_s_0_450 = 1.78e-05  mcm4m2_cc_w_2_400_s_0_450 = 9.79e-11  mcm4m2_cf_w_2_400_s_0_450 = 4.26e-12
+ mcm4m2_ca_w_2_400_s_0_600 = 1.78e-05  mcm4m2_cc_w_2_400_s_0_600 = 8.55e-11  mcm4m2_cf_w_2_400_s_0_600 = 5.47e-12
+ mcm4m2_ca_w_2_400_s_0_800 = 1.78e-05  mcm4m2_cc_w_2_400_s_0_800 = 7.31e-11  mcm4m2_cf_w_2_400_s_0_800 = 7.04e-12
+ mcm4m2_ca_w_2_400_s_1_000 = 1.78e-05  mcm4m2_cc_w_2_400_s_1_000 = 6.35e-11  mcm4m2_cf_w_2_400_s_1_000 = 8.55e-12
+ mcm4m2_ca_w_2_400_s_1_200 = 1.78e-05  mcm4m2_cc_w_2_400_s_1_200 = 5.64e-11  mcm4m2_cf_w_2_400_s_1_200 = 1.00e-11
+ mcm4m2_ca_w_2_400_s_2_100 = 1.78e-05  mcm4m2_cc_w_2_400_s_2_100 = 3.76e-11  mcm4m2_cf_w_2_400_s_2_100 = 1.58e-11
+ mcm4m2_ca_w_2_400_s_3_300 = 1.78e-05  mcm4m2_cc_w_2_400_s_3_300 = 2.55e-11  mcm4m2_cf_w_2_400_s_3_300 = 2.20e-11
+ mcm4m2_ca_w_2_400_s_9_000 = 1.78e-05  mcm4m2_cc_w_2_400_s_9_000 = 7.65e-12  mcm4m2_cf_w_2_400_s_9_000 = 3.60e-11
+ mcm4m3_ca_w_0_300_s_0_300 = 5.76e-05  mcm4m3_cc_w_0_300_s_0_300 = 8.23e-11  mcm4m3_cf_w_0_300_s_0_300 = 9.16e-12
+ mcm4m3_ca_w_0_300_s_0_360 = 5.76e-05  mcm4m3_cc_w_0_300_s_0_360 = 7.65e-11  mcm4m3_cf_w_0_300_s_0_360 = 1.06e-11
+ mcm4m3_ca_w_0_300_s_0_450 = 5.76e-05  mcm4m3_cc_w_0_300_s_0_450 = 6.85e-11  mcm4m3_cf_w_0_300_s_0_450 = 1.26e-11
+ mcm4m3_ca_w_0_300_s_0_600 = 5.76e-05  mcm4m3_cc_w_0_300_s_0_600 = 5.76e-11  mcm4m3_cf_w_0_300_s_0_600 = 1.58e-11
+ mcm4m3_ca_w_0_300_s_0_800 = 5.76e-05  mcm4m3_cc_w_0_300_s_0_800 = 4.72e-11  mcm4m3_cf_w_0_300_s_0_800 = 1.95e-11
+ mcm4m3_ca_w_0_300_s_1_000 = 5.76e-05  mcm4m3_cc_w_0_300_s_1_000 = 3.92e-11  mcm4m3_cf_w_0_300_s_1_000 = 2.28e-11
+ mcm4m3_ca_w_0_300_s_1_200 = 5.76e-05  mcm4m3_cc_w_0_300_s_1_200 = 3.31e-11  mcm4m3_cf_w_0_300_s_1_200 = 2.57e-11
+ mcm4m3_ca_w_0_300_s_2_100 = 5.76e-05  mcm4m3_cc_w_0_300_s_2_100 = 1.78e-11  mcm4m3_cf_w_0_300_s_2_100 = 3.57e-11
+ mcm4m3_ca_w_0_300_s_3_300 = 5.76e-05  mcm4m3_cc_w_0_300_s_3_300 = 1.02e-11  mcm4m3_cf_w_0_300_s_3_300 = 4.20e-11
+ mcm4m3_ca_w_0_300_s_9_000 = 5.76e-05  mcm4m3_cc_w_0_300_s_9_000 = 2.00e-12  mcm4m3_cf_w_0_300_s_9_000 = 4.98e-11
+ mcm4m3_ca_w_2_400_s_0_300 = 5.76e-05  mcm4m3_cc_w_2_400_s_0_300 = 1.01e-10  mcm4m3_cf_w_2_400_s_0_300 = 9.18e-12
+ mcm4m3_ca_w_2_400_s_0_360 = 5.76e-05  mcm4m3_cc_w_2_400_s_0_360 = 9.41e-11  mcm4m3_cf_w_2_400_s_0_360 = 1.06e-11
+ mcm4m3_ca_w_2_400_s_0_450 = 5.76e-05  mcm4m3_cc_w_2_400_s_0_450 = 8.51e-11  mcm4m3_cf_w_2_400_s_0_450 = 1.26e-11
+ mcm4m3_ca_w_2_400_s_0_600 = 5.76e-05  mcm4m3_cc_w_2_400_s_0_600 = 7.30e-11  mcm4m3_cf_w_2_400_s_0_600 = 1.58e-11
+ mcm4m3_ca_w_2_400_s_0_800 = 5.76e-05  mcm4m3_cc_w_2_400_s_0_800 = 6.08e-11  mcm4m3_cf_w_2_400_s_0_800 = 1.96e-11
+ mcm4m3_ca_w_2_400_s_1_000 = 5.76e-05  mcm4m3_cc_w_2_400_s_1_000 = 5.17e-11  mcm4m3_cf_w_2_400_s_1_000 = 2.29e-11
+ mcm4m3_ca_w_2_400_s_1_200 = 5.76e-05  mcm4m3_cc_w_2_400_s_1_200 = 4.47e-11  mcm4m3_cf_w_2_400_s_1_200 = 2.59e-11
+ mcm4m3_ca_w_2_400_s_2_100 = 5.76e-05  mcm4m3_cc_w_2_400_s_2_100 = 2.73e-11  mcm4m3_cf_w_2_400_s_2_100 = 3.58e-11
+ mcm4m3_ca_w_2_400_s_3_300 = 5.76e-05  mcm4m3_cc_w_2_400_s_3_300 = 1.68e-11  mcm4m3_cf_w_2_400_s_3_300 = 4.38e-11
+ mcm4m3_ca_w_2_400_s_9_000 = 5.76e-05  mcm4m3_cc_w_2_400_s_9_000 = 4.10e-12  mcm4m3_cf_w_2_400_s_9_000 = 5.57e-11
+ mcm5f_ca_w_1_600_s_1_600 = 5.56e-06  mcm5f_cc_w_1_600_s_1_600 = 6.47e-11  mcm5f_cf_w_1_600_s_1_600 = 4.59e-12
+ mcm5f_ca_w_1_600_s_1_700 = 5.56e-06  mcm5f_cc_w_1_600_s_1_700 = 6.19e-11  mcm5f_cf_w_1_600_s_1_700 = 4.85e-12
+ mcm5f_ca_w_1_600_s_1_900 = 5.56e-06  mcm5f_cc_w_1_600_s_1_900 = 5.72e-11  mcm5f_cf_w_1_600_s_1_900 = 5.36e-12
+ mcm5f_ca_w_1_600_s_2_000 = 5.56e-06  mcm5f_cc_w_1_600_s_2_000 = 5.52e-11  mcm5f_cf_w_1_600_s_2_000 = 5.61e-12
+ mcm5f_ca_w_1_600_s_2_400 = 5.56e-06  mcm5f_cc_w_1_600_s_2_400 = 4.85e-11  mcm5f_cf_w_1_600_s_2_400 = 6.60e-12
+ mcm5f_ca_w_1_600_s_2_800 = 5.56e-06  mcm5f_cc_w_1_600_s_2_800 = 4.33e-11  mcm5f_cf_w_1_600_s_2_800 = 7.57e-12
+ mcm5f_ca_w_1_600_s_3_200 = 5.56e-06  mcm5f_cc_w_1_600_s_3_200 = 3.93e-11  mcm5f_cf_w_1_600_s_3_200 = 8.50e-12
+ mcm5f_ca_w_1_600_s_4_800 = 5.56e-06  mcm5f_cc_w_1_600_s_4_800 = 2.87e-11  mcm5f_cf_w_1_600_s_4_800 = 1.20e-11
+ mcm5f_ca_w_1_600_s_10_000 = 5.56e-06  mcm5f_cc_w_1_600_s_10_000 = 1.42e-11  mcm5f_cf_w_1_600_s_10_000 = 2.02e-11
+ mcm5f_ca_w_1_600_s_12_000 = 5.56e-06  mcm5f_cc_w_1_600_s_12_000 = 1.14e-11  mcm5f_cf_w_1_600_s_12_000 = 2.23e-11
+ mcm5f_ca_w_4_000_s_1_600 = 5.56e-06  mcm5f_cc_w_4_000_s_1_600 = 7.24e-11  mcm5f_cf_w_4_000_s_1_600 = 4.60e-12
+ mcm5f_ca_w_4_000_s_1_700 = 5.56e-06  mcm5f_cc_w_4_000_s_1_700 = 6.93e-11  mcm5f_cf_w_4_000_s_1_700 = 4.86e-12
+ mcm5f_ca_w_4_000_s_1_900 = 5.56e-06  mcm5f_cc_w_4_000_s_1_900 = 6.42e-11  mcm5f_cf_w_4_000_s_1_900 = 5.37e-12
+ mcm5f_ca_w_4_000_s_2_000 = 5.56e-06  mcm5f_cc_w_4_000_s_2_000 = 6.19e-11  mcm5f_cf_w_4_000_s_2_000 = 5.62e-12
+ mcm5f_ca_w_4_000_s_2_400 = 5.56e-06  mcm5f_cc_w_4_000_s_2_400 = 5.46e-11  mcm5f_cf_w_4_000_s_2_400 = 6.61e-12
+ mcm5f_ca_w_4_000_s_2_800 = 5.56e-06  mcm5f_cc_w_4_000_s_2_800 = 4.91e-11  mcm5f_cf_w_4_000_s_2_800 = 7.59e-12
+ mcm5f_ca_w_4_000_s_3_200 = 5.56e-06  mcm5f_cc_w_4_000_s_3_200 = 4.47e-11  mcm5f_cf_w_4_000_s_3_200 = 8.53e-12
+ mcm5f_ca_w_4_000_s_4_800 = 5.56e-06  mcm5f_cc_w_4_000_s_4_800 = 3.30e-11  mcm5f_cf_w_4_000_s_4_800 = 1.20e-11
+ mcm5f_ca_w_4_000_s_10_000 = 5.56e-06  mcm5f_cc_w_4_000_s_10_000 = 1.70e-11  mcm5f_cf_w_4_000_s_10_000 = 2.06e-11
+ mcm5f_ca_w_4_000_s_12_000 = 5.56e-06  mcm5f_cc_w_4_000_s_12_000 = 1.39e-11  mcm5f_cf_w_4_000_s_12_000 = 2.29e-11
+ mcm5d_ca_w_1_600_s_1_600 = 5.96e-06  mcm5d_cc_w_1_600_s_1_600 = 6.42e-11  mcm5d_cf_w_1_600_s_1_600 = 4.91e-12
+ mcm5d_ca_w_1_600_s_1_700 = 5.96e-06  mcm5d_cc_w_1_600_s_1_700 = 6.15e-11  mcm5d_cf_w_1_600_s_1_700 = 5.18e-12
+ mcm5d_ca_w_1_600_s_1_900 = 5.96e-06  mcm5d_cc_w_1_600_s_1_900 = 5.67e-11  mcm5d_cf_w_1_600_s_1_900 = 5.73e-12
+ mcm5d_ca_w_1_600_s_2_000 = 5.96e-06  mcm5d_cc_w_1_600_s_2_000 = 5.47e-11  mcm5d_cf_w_1_600_s_2_000 = 5.99e-12
+ mcm5d_ca_w_1_600_s_2_400 = 5.96e-06  mcm5d_cc_w_1_600_s_2_400 = 4.79e-11  mcm5d_cf_w_1_600_s_2_400 = 7.04e-12
+ mcm5d_ca_w_1_600_s_2_800 = 5.96e-06  mcm5d_cc_w_1_600_s_2_800 = 4.28e-11  mcm5d_cf_w_1_600_s_2_800 = 8.07e-12
+ mcm5d_ca_w_1_600_s_3_200 = 5.96e-06  mcm5d_cc_w_1_600_s_3_200 = 3.88e-11  mcm5d_cf_w_1_600_s_3_200 = 9.06e-12
+ mcm5d_ca_w_1_600_s_4_800 = 5.96e-06  mcm5d_cc_w_1_600_s_4_800 = 2.81e-11  mcm5d_cf_w_1_600_s_4_800 = 1.27e-11
+ mcm5d_ca_w_1_600_s_10_000 = 5.96e-06  mcm5d_cc_w_1_600_s_10_000 = 1.36e-11  mcm5d_cf_w_1_600_s_10_000 = 2.12e-11
+ mcm5d_ca_w_1_600_s_12_000 = 5.96e-06  mcm5d_cc_w_1_600_s_12_000 = 1.09e-11  mcm5d_cf_w_1_600_s_12_000 = 2.33e-11
+ mcm5d_ca_w_4_000_s_1_600 = 5.96e-06  mcm5d_cc_w_4_000_s_1_600 = 7.18e-11  mcm5d_cf_w_4_000_s_1_600 = 4.92e-12
+ mcm5d_ca_w_4_000_s_1_700 = 5.96e-06  mcm5d_cc_w_4_000_s_1_700 = 6.87e-11  mcm5d_cf_w_4_000_s_1_700 = 5.20e-12
+ mcm5d_ca_w_4_000_s_1_900 = 5.96e-06  mcm5d_cc_w_4_000_s_1_900 = 6.35e-11  mcm5d_cf_w_4_000_s_1_900 = 5.74e-12
+ mcm5d_ca_w_4_000_s_2_000 = 5.96e-06  mcm5d_cc_w_4_000_s_2_000 = 6.13e-11  mcm5d_cf_w_4_000_s_2_000 = 6.00e-12
+ mcm5d_ca_w_4_000_s_2_400 = 5.96e-06  mcm5d_cc_w_4_000_s_2_400 = 5.39e-11  mcm5d_cf_w_4_000_s_2_400 = 7.05e-12
+ mcm5d_ca_w_4_000_s_2_800 = 5.96e-06  mcm5d_cc_w_4_000_s_2_800 = 4.84e-11  mcm5d_cf_w_4_000_s_2_800 = 8.09e-12
+ mcm5d_ca_w_4_000_s_3_200 = 5.96e-06  mcm5d_cc_w_4_000_s_3_200 = 4.40e-11  mcm5d_cf_w_4_000_s_3_200 = 9.09e-12
+ mcm5d_ca_w_4_000_s_4_800 = 5.96e-06  mcm5d_cc_w_4_000_s_4_800 = 3.23e-11  mcm5d_cf_w_4_000_s_4_800 = 1.28e-11
+ mcm5d_ca_w_4_000_s_10_000 = 5.96e-06  mcm5d_cc_w_4_000_s_10_000 = 1.64e-11  mcm5d_cf_w_4_000_s_10_000 = 2.17e-11
+ mcm5d_ca_w_4_000_s_12_000 = 5.96e-06  mcm5d_cc_w_4_000_s_12_000 = 1.34e-11  mcm5d_cf_w_4_000_s_12_000 = 2.40e-11
+ mcm5p1_ca_w_1_600_s_1_600 = 6.20e-06  mcm5p1_cc_w_1_600_s_1_600 = 6.41e-11  mcm5p1_cf_w_1_600_s_1_600 = 5.11e-12
+ mcm5p1_ca_w_1_600_s_1_700 = 6.20e-06  mcm5p1_cc_w_1_600_s_1_700 = 6.13e-11  mcm5p1_cf_w_1_600_s_1_700 = 5.39e-12
+ mcm5p1_ca_w_1_600_s_1_900 = 6.20e-06  mcm5p1_cc_w_1_600_s_1_900 = 5.64e-11  mcm5p1_cf_w_1_600_s_1_900 = 5.96e-12
+ mcm5p1_ca_w_1_600_s_2_000 = 6.20e-06  mcm5p1_cc_w_1_600_s_2_000 = 5.44e-11  mcm5p1_cf_w_1_600_s_2_000 = 6.23e-12
+ mcm5p1_ca_w_1_600_s_2_400 = 6.20e-06  mcm5p1_cc_w_1_600_s_2_400 = 4.76e-11  mcm5p1_cf_w_1_600_s_2_400 = 7.32e-12
+ mcm5p1_ca_w_1_600_s_2_800 = 6.20e-06  mcm5p1_cc_w_1_600_s_2_800 = 4.24e-11  mcm5p1_cf_w_1_600_s_2_800 = 8.38e-12
+ mcm5p1_ca_w_1_600_s_3_200 = 6.20e-06  mcm5p1_cc_w_1_600_s_3_200 = 3.84e-11  mcm5p1_cf_w_1_600_s_3_200 = 9.41e-12
+ mcm5p1_ca_w_1_600_s_4_800 = 6.20e-06  mcm5p1_cc_w_1_600_s_4_800 = 2.77e-11  mcm5p1_cf_w_1_600_s_4_800 = 1.31e-11
+ mcm5p1_ca_w_1_600_s_10_000 = 6.20e-06  mcm5p1_cc_w_1_600_s_10_000 = 1.33e-11  mcm5p1_cf_w_1_600_s_10_000 = 2.18e-11
+ mcm5p1_ca_w_1_600_s_12_000 = 6.20e-06  mcm5p1_cc_w_1_600_s_12_000 = 1.06e-11  mcm5p1_cf_w_1_600_s_12_000 = 2.39e-11
+ mcm5p1_ca_w_4_000_s_1_600 = 6.20e-06  mcm5p1_cc_w_4_000_s_1_600 = 7.14e-11  mcm5p1_cf_w_4_000_s_1_600 = 5.12e-12
+ mcm5p1_ca_w_4_000_s_1_700 = 6.20e-06  mcm5p1_cc_w_4_000_s_1_700 = 6.83e-11  mcm5p1_cf_w_4_000_s_1_700 = 5.41e-12
+ mcm5p1_ca_w_4_000_s_1_900 = 6.20e-06  mcm5p1_cc_w_4_000_s_1_900 = 6.31e-11  mcm5p1_cf_w_4_000_s_1_900 = 5.97e-12
+ mcm5p1_ca_w_4_000_s_2_000 = 6.20e-06  mcm5p1_cc_w_4_000_s_2_000 = 6.09e-11  mcm5p1_cf_w_4_000_s_2_000 = 6.24e-12
+ mcm5p1_ca_w_4_000_s_2_400 = 6.20e-06  mcm5p1_cc_w_4_000_s_2_400 = 5.36e-11  mcm5p1_cf_w_4_000_s_2_400 = 7.33e-12
+ mcm5p1_ca_w_4_000_s_2_800 = 6.20e-06  mcm5p1_cc_w_4_000_s_2_800 = 4.80e-11  mcm5p1_cf_w_4_000_s_2_800 = 8.40e-12
+ mcm5p1_ca_w_4_000_s_3_200 = 6.20e-06  mcm5p1_cc_w_4_000_s_3_200 = 4.35e-11  mcm5p1_cf_w_4_000_s_3_200 = 9.44e-12
+ mcm5p1_ca_w_4_000_s_4_800 = 6.20e-06  mcm5p1_cc_w_4_000_s_4_800 = 3.19e-11  mcm5p1_cf_w_4_000_s_4_800 = 1.32e-11
+ mcm5p1_ca_w_4_000_s_10_000 = 6.20e-06  mcm5p1_cc_w_4_000_s_10_000 = 1.61e-11  mcm5p1_cf_w_4_000_s_10_000 = 2.23e-11
+ mcm5p1_ca_w_4_000_s_12_000 = 6.20e-06  mcm5p1_cc_w_4_000_s_12_000 = 1.30e-11  mcm5p1_cf_w_4_000_s_12_000 = 2.46e-11
+ mcm5l1_ca_w_1_600_s_1_600 = 6.97e-06  mcm5l1_cc_w_1_600_s_1_600 = 6.32e-11  mcm5l1_cf_w_1_600_s_1_600 = 5.71e-12
+ mcm5l1_ca_w_1_600_s_1_700 = 6.97e-06  mcm5l1_cc_w_1_600_s_1_700 = 6.05e-11  mcm5l1_cf_w_1_600_s_1_700 = 6.02e-12
+ mcm5l1_ca_w_1_600_s_1_900 = 6.97e-06  mcm5l1_cc_w_1_600_s_1_900 = 5.56e-11  mcm5l1_cf_w_1_600_s_1_900 = 6.65e-12
+ mcm5l1_ca_w_1_600_s_2_000 = 6.97e-06  mcm5l1_cc_w_1_600_s_2_000 = 5.35e-11  mcm5l1_cf_w_1_600_s_2_000 = 6.96e-12
+ mcm5l1_ca_w_1_600_s_2_400 = 6.97e-06  mcm5l1_cc_w_1_600_s_2_400 = 4.67e-11  mcm5l1_cf_w_1_600_s_2_400 = 8.16e-12
+ mcm5l1_ca_w_1_600_s_2_800 = 6.97e-06  mcm5l1_cc_w_1_600_s_2_800 = 4.15e-11  mcm5l1_cf_w_1_600_s_2_800 = 9.33e-12
+ mcm5l1_ca_w_1_600_s_3_200 = 6.97e-06  mcm5l1_cc_w_1_600_s_3_200 = 3.74e-11  mcm5l1_cf_w_1_600_s_3_200 = 1.05e-11
+ mcm5l1_ca_w_1_600_s_4_800 = 6.97e-06  mcm5l1_cc_w_1_600_s_4_800 = 2.67e-11  mcm5l1_cf_w_1_600_s_4_800 = 1.45e-11
+ mcm5l1_ca_w_1_600_s_10_000 = 6.97e-06  mcm5l1_cc_w_1_600_s_10_000 = 1.24e-11  mcm5l1_cf_w_1_600_s_10_000 = 2.35e-11
+ mcm5l1_ca_w_1_600_s_12_000 = 6.97e-06  mcm5l1_cc_w_1_600_s_12_000 = 9.77e-12  mcm5l1_cf_w_1_600_s_12_000 = 2.57e-11
+ mcm5l1_ca_w_4_000_s_1_600 = 6.97e-06  mcm5l1_cc_w_4_000_s_1_600 = 7.02e-11  mcm5l1_cf_w_4_000_s_1_600 = 5.71e-12
+ mcm5l1_ca_w_4_000_s_1_700 = 6.97e-06  mcm5l1_cc_w_4_000_s_1_700 = 6.72e-11  mcm5l1_cf_w_4_000_s_1_700 = 6.04e-12
+ mcm5l1_ca_w_4_000_s_1_900 = 6.97e-06  mcm5l1_cc_w_4_000_s_1_900 = 6.20e-11  mcm5l1_cf_w_4_000_s_1_900 = 6.66e-12
+ mcm5l1_ca_w_4_000_s_2_000 = 6.97e-06  mcm5l1_cc_w_4_000_s_2_000 = 5.97e-11  mcm5l1_cf_w_4_000_s_2_000 = 6.97e-12
+ mcm5l1_ca_w_4_000_s_2_400 = 6.97e-06  mcm5l1_cc_w_4_000_s_2_400 = 5.24e-11  mcm5l1_cf_w_4_000_s_2_400 = 8.17e-12
+ mcm5l1_ca_w_4_000_s_2_800 = 6.97e-06  mcm5l1_cc_w_4_000_s_2_800 = 4.68e-11  mcm5l1_cf_w_4_000_s_2_800 = 9.35e-12
+ mcm5l1_ca_w_4_000_s_3_200 = 6.97e-06  mcm5l1_cc_w_4_000_s_3_200 = 4.24e-11  mcm5l1_cf_w_4_000_s_3_200 = 1.05e-11
+ mcm5l1_ca_w_4_000_s_4_800 = 6.97e-06  mcm5l1_cc_w_4_000_s_4_800 = 3.07e-11  mcm5l1_cf_w_4_000_s_4_800 = 1.46e-11
+ mcm5l1_ca_w_4_000_s_10_000 = 6.97e-06  mcm5l1_cc_w_4_000_s_10_000 = 1.51e-11  mcm5l1_cf_w_4_000_s_10_000 = 2.41e-11
+ mcm5l1_ca_w_4_000_s_12_000 = 6.97e-06  mcm5l1_cc_w_4_000_s_12_000 = 1.21e-11  mcm5l1_cf_w_4_000_s_12_000 = 2.64e-11
+ mcm5m1_ca_w_1_600_s_1_600 = 8.26e-06  mcm5m1_cc_w_1_600_s_1_600 = 6.19e-11  mcm5m1_cf_w_1_600_s_1_600 = 6.71e-12
+ mcm5m1_ca_w_1_600_s_1_700 = 8.26e-06  mcm5m1_cc_w_1_600_s_1_700 = 5.91e-11  mcm5m1_cf_w_1_600_s_1_700 = 7.07e-12
+ mcm5m1_ca_w_1_600_s_1_900 = 8.26e-06  mcm5m1_cc_w_1_600_s_1_900 = 5.42e-11  mcm5m1_cf_w_1_600_s_1_900 = 7.80e-12
+ mcm5m1_ca_w_1_600_s_2_000 = 8.26e-06  mcm5m1_cc_w_1_600_s_2_000 = 5.21e-11  mcm5m1_cf_w_1_600_s_2_000 = 8.16e-12
+ mcm5m1_ca_w_1_600_s_2_400 = 8.26e-06  mcm5m1_cc_w_1_600_s_2_400 = 4.53e-11  mcm5m1_cf_w_1_600_s_2_400 = 9.55e-12
+ mcm5m1_ca_w_1_600_s_2_800 = 8.26e-06  mcm5m1_cc_w_1_600_s_2_800 = 4.00e-11  mcm5m1_cf_w_1_600_s_2_800 = 1.09e-11
+ mcm5m1_ca_w_1_600_s_3_200 = 8.26e-06  mcm5m1_cc_w_1_600_s_3_200 = 3.59e-11  mcm5m1_cf_w_1_600_s_3_200 = 1.22e-11
+ mcm5m1_ca_w_1_600_s_4_800 = 8.26e-06  mcm5m1_cc_w_1_600_s_4_800 = 2.51e-11  mcm5m1_cf_w_1_600_s_4_800 = 1.67e-11
+ mcm5m1_ca_w_1_600_s_10_000 = 8.26e-06  mcm5m1_cc_w_1_600_s_10_000 = 1.11e-11  mcm5m1_cf_w_1_600_s_10_000 = 2.62e-11
+ mcm5m1_ca_w_1_600_s_12_000 = 8.26e-06  mcm5m1_cc_w_1_600_s_12_000 = 8.66e-12  mcm5m1_cf_w_1_600_s_12_000 = 2.83e-11
+ mcm5m1_ca_w_4_000_s_1_600 = 8.26e-06  mcm5m1_cc_w_4_000_s_1_600 = 6.85e-11  mcm5m1_cf_w_4_000_s_1_600 = 6.71e-12
+ mcm5m1_ca_w_4_000_s_1_700 = 8.26e-06  mcm5m1_cc_w_4_000_s_1_700 = 6.55e-11  mcm5m1_cf_w_4_000_s_1_700 = 7.10e-12
+ mcm5m1_ca_w_4_000_s_1_900 = 8.26e-06  mcm5m1_cc_w_4_000_s_1_900 = 6.04e-11  mcm5m1_cf_w_4_000_s_1_900 = 7.82e-12
+ mcm5m1_ca_w_4_000_s_2_000 = 8.26e-06  mcm5m1_cc_w_4_000_s_2_000 = 5.80e-11  mcm5m1_cf_w_4_000_s_2_000 = 8.17e-12
+ mcm5m1_ca_w_4_000_s_2_400 = 8.26e-06  mcm5m1_cc_w_4_000_s_2_400 = 5.07e-11  mcm5m1_cf_w_4_000_s_2_400 = 9.56e-12
+ mcm5m1_ca_w_4_000_s_2_800 = 8.26e-06  mcm5m1_cc_w_4_000_s_2_800 = 4.51e-11  mcm5m1_cf_w_4_000_s_2_800 = 1.09e-11
+ mcm5m1_ca_w_4_000_s_3_200 = 8.26e-06  mcm5m1_cc_w_4_000_s_3_200 = 4.07e-11  mcm5m1_cf_w_4_000_s_3_200 = 1.22e-11
+ mcm5m1_ca_w_4_000_s_4_800 = 8.26e-06  mcm5m1_cc_w_4_000_s_4_800 = 2.90e-11  mcm5m1_cf_w_4_000_s_4_800 = 1.68e-11
+ mcm5m1_ca_w_4_000_s_10_000 = 8.26e-06  mcm5m1_cc_w_4_000_s_10_000 = 1.37e-11  mcm5m1_cf_w_4_000_s_10_000 = 2.68e-11
+ mcm5m1_ca_w_4_000_s_12_000 = 8.26e-06  mcm5m1_cc_w_4_000_s_12_000 = 1.09e-11  mcm5m1_cf_w_4_000_s_12_000 = 2.92e-11
+ mcm5m2_ca_w_1_600_s_1_600 = 1.01e-05  mcm5m2_cc_w_1_600_s_1_600 = 6.03e-11  mcm5m2_cf_w_1_600_s_1_600 = 8.11e-12
+ mcm5m2_ca_w_1_600_s_1_700 = 1.01e-05  mcm5m2_cc_w_1_600_s_1_700 = 5.74e-11  mcm5m2_cf_w_1_600_s_1_700 = 8.54e-12
+ mcm5m2_ca_w_1_600_s_1_900 = 1.01e-05  mcm5m2_cc_w_1_600_s_1_900 = 5.25e-11  mcm5m2_cf_w_1_600_s_1_900 = 9.40e-12
+ mcm5m2_ca_w_1_600_s_2_000 = 1.01e-05  mcm5m2_cc_w_1_600_s_2_000 = 5.04e-11  mcm5m2_cf_w_1_600_s_2_000 = 9.82e-12
+ mcm5m2_ca_w_1_600_s_2_400 = 1.01e-05  mcm5m2_cc_w_1_600_s_2_400 = 4.35e-11  mcm5m2_cf_w_1_600_s_2_400 = 1.15e-11
+ mcm5m2_ca_w_1_600_s_2_800 = 1.01e-05  mcm5m2_cc_w_1_600_s_2_800 = 3.82e-11  mcm5m2_cf_w_1_600_s_2_800 = 1.30e-11
+ mcm5m2_ca_w_1_600_s_3_200 = 1.01e-05  mcm5m2_cc_w_1_600_s_3_200 = 3.40e-11  mcm5m2_cf_w_1_600_s_3_200 = 1.45e-11
+ mcm5m2_ca_w_1_600_s_4_800 = 1.01e-05  mcm5m2_cc_w_1_600_s_4_800 = 2.33e-11  mcm5m2_cf_w_1_600_s_4_800 = 1.96e-11
+ mcm5m2_ca_w_1_600_s_10_000 = 1.01e-05  mcm5m2_cc_w_1_600_s_10_000 = 9.71e-12  mcm5m2_cf_w_1_600_s_10_000 = 2.95e-11
+ mcm5m2_ca_w_1_600_s_12_000 = 1.01e-05  mcm5m2_cc_w_1_600_s_12_000 = 7.44e-12  mcm5m2_cf_w_1_600_s_12_000 = 3.15e-11
+ mcm5m2_ca_w_4_000_s_1_600 = 1.01e-05  mcm5m2_cc_w_4_000_s_1_600 = 6.64e-11  mcm5m2_cf_w_4_000_s_1_600 = 8.11e-12
+ mcm5m2_ca_w_4_000_s_1_700 = 1.01e-05  mcm5m2_cc_w_4_000_s_1_700 = 6.34e-11  mcm5m2_cf_w_4_000_s_1_700 = 8.55e-12
+ mcm5m2_ca_w_4_000_s_1_900 = 1.01e-05  mcm5m2_cc_w_4_000_s_1_900 = 5.83e-11  mcm5m2_cf_w_4_000_s_1_900 = 9.41e-12
+ mcm5m2_ca_w_4_000_s_2_000 = 1.01e-05  mcm5m2_cc_w_4_000_s_2_000 = 5.60e-11  mcm5m2_cf_w_4_000_s_2_000 = 9.84e-12
+ mcm5m2_ca_w_4_000_s_2_400 = 1.01e-05  mcm5m2_cc_w_4_000_s_2_400 = 4.86e-11  mcm5m2_cf_w_4_000_s_2_400 = 1.15e-11
+ mcm5m2_ca_w_4_000_s_2_800 = 1.01e-05  mcm5m2_cc_w_4_000_s_2_800 = 4.30e-11  mcm5m2_cf_w_4_000_s_2_800 = 1.30e-11
+ mcm5m2_ca_w_4_000_s_3_200 = 1.01e-05  mcm5m2_cc_w_4_000_s_3_200 = 3.86e-11  mcm5m2_cf_w_4_000_s_3_200 = 1.45e-11
+ mcm5m2_ca_w_4_000_s_4_800 = 1.01e-05  mcm5m2_cc_w_4_000_s_4_800 = 2.71e-11  mcm5m2_cf_w_4_000_s_4_800 = 1.97e-11
+ mcm5m2_ca_w_4_000_s_10_000 = 1.01e-05  mcm5m2_cc_w_4_000_s_10_000 = 1.22e-11  mcm5m2_cf_w_4_000_s_10_000 = 3.02e-11
+ mcm5m2_ca_w_4_000_s_12_000 = 1.01e-05  mcm5m2_cc_w_4_000_s_12_000 = 9.60e-12  mcm5m2_cf_w_4_000_s_12_000 = 3.24e-11
+ mcm5m3_ca_w_1_600_s_1_600 = 1.67e-05  mcm5m3_cc_w_1_600_s_1_600 = 5.54e-11  mcm5m3_cf_w_1_600_s_1_600 = 1.28e-11
+ mcm5m3_ca_w_1_600_s_1_700 = 1.67e-05  mcm5m3_cc_w_1_600_s_1_700 = 5.26e-11  mcm5m3_cf_w_1_600_s_1_700 = 1.35e-11
+ mcm5m3_ca_w_1_600_s_1_900 = 1.67e-05  mcm5m3_cc_w_1_600_s_1_900 = 4.76e-11  mcm5m3_cf_w_1_600_s_1_900 = 1.48e-11
+ mcm5m3_ca_w_1_600_s_2_000 = 1.67e-05  mcm5m3_cc_w_1_600_s_2_000 = 4.55e-11  mcm5m3_cf_w_1_600_s_2_000 = 1.54e-11
+ mcm5m3_ca_w_1_600_s_2_400 = 1.67e-05  mcm5m3_cc_w_1_600_s_2_400 = 3.85e-11  mcm5m3_cf_w_1_600_s_2_400 = 1.77e-11
+ mcm5m3_ca_w_1_600_s_2_800 = 1.67e-05  mcm5m3_cc_w_1_600_s_2_800 = 3.33e-11  mcm5m3_cf_w_1_600_s_2_800 = 1.99e-11
+ mcm5m3_ca_w_1_600_s_3_200 = 1.67e-05  mcm5m3_cc_w_1_600_s_3_200 = 2.92e-11  mcm5m3_cf_w_1_600_s_3_200 = 2.19e-11
+ mcm5m3_ca_w_1_600_s_4_800 = 1.67e-05  mcm5m3_cc_w_1_600_s_4_800 = 1.88e-11  mcm5m3_cf_w_1_600_s_4_800 = 2.82e-11
+ mcm5m3_ca_w_1_600_s_10_000 = 1.67e-05  mcm5m3_cc_w_1_600_s_10_000 = 6.95e-12  mcm5m3_cf_w_1_600_s_10_000 = 3.81e-11
+ mcm5m3_ca_w_1_600_s_12_000 = 1.67e-05  mcm5m3_cc_w_1_600_s_12_000 = 5.20e-12  mcm5m3_cf_w_1_600_s_12_000 = 3.97e-11
+ mcm5m3_ca_w_4_000_s_1_600 = 1.67e-05  mcm5m3_cc_w_4_000_s_1_600 = 6.09e-11  mcm5m3_cf_w_4_000_s_1_600 = 1.28e-11
+ mcm5m3_ca_w_4_000_s_1_700 = 1.67e-05  mcm5m3_cc_w_4_000_s_1_700 = 5.81e-11  mcm5m3_cf_w_4_000_s_1_700 = 1.35e-11
+ mcm5m3_ca_w_4_000_s_1_900 = 1.67e-05  mcm5m3_cc_w_4_000_s_1_900 = 5.29e-11  mcm5m3_cf_w_4_000_s_1_900 = 1.48e-11
+ mcm5m3_ca_w_4_000_s_2_000 = 1.67e-05  mcm5m3_cc_w_4_000_s_2_000 = 5.07e-11  mcm5m3_cf_w_4_000_s_2_000 = 1.54e-11
+ mcm5m3_ca_w_4_000_s_2_400 = 1.67e-05  mcm5m3_cc_w_4_000_s_2_400 = 4.33e-11  mcm5m3_cf_w_4_000_s_2_400 = 1.77e-11
+ mcm5m3_ca_w_4_000_s_2_800 = 1.67e-05  mcm5m3_cc_w_4_000_s_2_800 = 3.78e-11  mcm5m3_cf_w_4_000_s_2_800 = 1.99e-11
+ mcm5m3_ca_w_4_000_s_3_200 = 1.67e-05  mcm5m3_cc_w_4_000_s_3_200 = 3.35e-11  mcm5m3_cf_w_4_000_s_3_200 = 2.19e-11
+ mcm5m3_ca_w_4_000_s_4_800 = 1.67e-05  mcm5m3_cc_w_4_000_s_4_800 = 2.24e-11  mcm5m3_cf_w_4_000_s_4_800 = 2.84e-11
+ mcm5m3_ca_w_4_000_s_10_000 = 1.67e-05  mcm5m3_cc_w_4_000_s_10_000 = 9.25e-12  mcm5m3_cf_w_4_000_s_10_000 = 3.90e-11
+ mcm5m3_ca_w_4_000_s_12_000 = 1.67e-05  mcm5m3_cc_w_4_000_s_12_000 = 7.15e-12  mcm5m3_cf_w_4_000_s_12_000 = 4.09e-11
+ mcm5m4_ca_w_1_600_s_1_600 = 4.87e-05  mcm5m4_cc_w_1_600_s_1_600 = 4.44e-11  mcm5m4_cf_w_1_600_s_1_600 = 3.09e-11
+ mcm5m4_ca_w_1_600_s_1_700 = 4.87e-05  mcm5m4_cc_w_1_600_s_1_700 = 4.16e-11  mcm5m4_cf_w_1_600_s_1_700 = 3.21e-11
+ mcm5m4_ca_w_1_600_s_1_900 = 4.87e-05  mcm5m4_cc_w_1_600_s_1_900 = 3.70e-11  mcm5m4_cf_w_1_600_s_1_900 = 3.44e-11
+ mcm5m4_ca_w_1_600_s_2_000 = 4.87e-05  mcm5m4_cc_w_1_600_s_2_000 = 3.50e-11  mcm5m4_cf_w_1_600_s_2_000 = 3.54e-11
+ mcm5m4_ca_w_1_600_s_2_400 = 4.87e-05  mcm5m4_cc_w_1_600_s_2_400 = 2.85e-11  mcm5m4_cf_w_1_600_s_2_400 = 3.91e-11
+ mcm5m4_ca_w_1_600_s_2_800 = 4.87e-05  mcm5m4_cc_w_1_600_s_2_800 = 2.38e-11  mcm5m4_cf_w_1_600_s_2_800 = 4.22e-11
+ mcm5m4_ca_w_1_600_s_3_200 = 4.87e-05  mcm5m4_cc_w_1_600_s_3_200 = 2.02e-11  mcm5m4_cf_w_1_600_s_3_200 = 4.47e-11
+ mcm5m4_ca_w_1_600_s_4_800 = 4.87e-05  mcm5m4_cc_w_1_600_s_4_800 = 1.19e-11  mcm5m4_cf_w_1_600_s_4_800 = 5.15e-11
+ mcm5m4_ca_w_1_600_s_10_000 = 4.87e-05  mcm5m4_cc_w_1_600_s_10_000 = 4.00e-12  mcm5m4_cf_w_1_600_s_10_000 = 5.89e-11
+ mcm5m4_ca_w_1_600_s_12_000 = 4.87e-05  mcm5m4_cc_w_1_600_s_12_000 = 2.95e-12  mcm5m4_cf_w_1_600_s_12_000 = 5.99e-11
+ mcm5m4_ca_w_4_000_s_1_600 = 4.87e-05  mcm5m4_cc_w_4_000_s_1_600 = 4.98e-11  mcm5m4_cf_w_4_000_s_1_600 = 3.09e-11
+ mcm5m4_ca_w_4_000_s_1_700 = 4.87e-05  mcm5m4_cc_w_4_000_s_1_700 = 4.70e-11  mcm5m4_cf_w_4_000_s_1_700 = 3.21e-11
+ mcm5m4_ca_w_4_000_s_1_900 = 4.87e-05  mcm5m4_cc_w_4_000_s_1_900 = 4.21e-11  mcm5m4_cf_w_4_000_s_1_900 = 3.44e-11
+ mcm5m4_ca_w_4_000_s_2_000 = 4.87e-05  mcm5m4_cc_w_4_000_s_2_000 = 4.00e-11  mcm5m4_cf_w_4_000_s_2_000 = 3.54e-11
+ mcm5m4_ca_w_4_000_s_2_400 = 4.87e-05  mcm5m4_cc_w_4_000_s_2_400 = 3.32e-11  mcm5m4_cf_w_4_000_s_2_400 = 3.91e-11
+ mcm5m4_ca_w_4_000_s_2_800 = 4.87e-05  mcm5m4_cc_w_4_000_s_2_800 = 2.83e-11  mcm5m4_cf_w_4_000_s_2_800 = 4.23e-11
+ mcm5m4_ca_w_4_000_s_3_200 = 4.87e-05  mcm5m4_cc_w_4_000_s_3_200 = 2.45e-11  mcm5m4_cf_w_4_000_s_3_200 = 4.49e-11
+ mcm5m4_ca_w_4_000_s_4_800 = 4.87e-05  mcm5m4_cc_w_4_000_s_4_800 = 1.55e-11  mcm5m4_cf_w_4_000_s_4_800 = 5.19e-11
+ mcm5m4_ca_w_4_000_s_10_000 = 4.87e-05  mcm5m4_cc_w_4_000_s_10_000 = 6.05e-12  mcm5m4_cf_w_4_000_s_10_000 = 6.06e-11
+ mcm5m4_ca_w_4_000_s_12_000 = 4.87e-05  mcm5m4_cc_w_4_000_s_12_000 = 4.70e-12  mcm5m4_cf_w_4_000_s_12_000 = 6.20e-11
+ mcrdlf_ca_w_10_000_s_5_000 = 2.15e-06  mcrdlf_cc_w_10_000_s_5_000 = 4.11e-11  mcrdlf_cf_w_10_000_s_5_000 = 5.98e-12
+ mcrdlf_ca_w_10_000_s_8_000 = 2.15e-06  mcrdlf_cc_w_10_000_s_8_000 = 3.16e-11  mcrdlf_cf_w_10_000_s_8_000 = 8.54e-12
+ mcrdlf_ca_w_10_000_s_10_000 = 2.15e-06  mcrdlf_cc_w_10_000_s_10_000 = 2.75e-11  mcrdlf_cf_w_10_000_s_10_000 = 1.01e-11
+ mcrdlf_ca_w_10_000_s_12_000 = 2.15e-06  mcrdlf_cc_w_10_000_s_12_000 = 2.44e-11  mcrdlf_cf_w_10_000_s_12_000 = 1.15e-11
+ mcrdlf_ca_w_10_000_s_30_000 = 2.15e-06  mcrdlf_cc_w_10_000_s_30_000 = 1.12e-11  mcrdlf_cf_w_10_000_s_30_000 = 2.04e-11
+ mcrdlf_ca_w_40_000_s_5_000 = 2.15e-06  mcrdlf_cc_w_40_000_s_5_000 = 5.25e-11  mcrdlf_cf_w_40_000_s_5_000 = 6.05e-12
+ mcrdlf_ca_w_40_000_s_8_000 = 2.15e-06  mcrdlf_cc_w_40_000_s_8_000 = 4.20e-11  mcrdlf_cf_w_40_000_s_8_000 = 8.63e-12
+ mcrdlf_ca_w_40_000_s_10_000 = 2.15e-06  mcrdlf_cc_w_40_000_s_10_000 = 3.74e-11  mcrdlf_cf_w_40_000_s_10_000 = 1.02e-11
+ mcrdlf_ca_w_40_000_s_12_000 = 2.15e-06  mcrdlf_cc_w_40_000_s_12_000 = 3.39e-11  mcrdlf_cf_w_40_000_s_12_000 = 1.17e-11
+ mcrdlf_ca_w_40_000_s_30_000 = 2.15e-06  mcrdlf_cc_w_40_000_s_30_000 = 1.84e-11  mcrdlf_cf_w_40_000_s_30_000 = 2.12e-11
+ mcrdld_ca_w_10_000_s_5_000 = 2.21e-06  mcrdld_cc_w_10_000_s_5_000 = 4.09e-11  mcrdld_cf_w_10_000_s_5_000 = 6.11e-12
+ mcrdld_ca_w_10_000_s_8_000 = 2.21e-06  mcrdld_cc_w_10_000_s_8_000 = 3.14e-11  mcrdld_cf_w_10_000_s_8_000 = 8.74e-12
+ mcrdld_ca_w_10_000_s_10_000 = 2.21e-06  mcrdld_cc_w_10_000_s_10_000 = 2.73e-11  mcrdld_cf_w_10_000_s_10_000 = 1.03e-11
+ mcrdld_ca_w_10_000_s_12_000 = 2.21e-06  mcrdld_cc_w_10_000_s_12_000 = 2.41e-11  mcrdld_cf_w_10_000_s_12_000 = 1.18e-11
+ mcrdld_ca_w_10_000_s_30_000 = 2.21e-06  mcrdld_cc_w_10_000_s_30_000 = 1.10e-11  mcrdld_cf_w_10_000_s_30_000 = 2.07e-11
+ mcrdld_ca_w_40_000_s_5_000 = 2.21e-06  mcrdld_cc_w_40_000_s_5_000 = 5.23e-11  mcrdld_cf_w_40_000_s_5_000 = 6.19e-12
+ mcrdld_ca_w_40_000_s_8_000 = 2.21e-06  mcrdld_cc_w_40_000_s_8_000 = 4.18e-11  mcrdld_cf_w_40_000_s_8_000 = 8.83e-12
+ mcrdld_ca_w_40_000_s_10_000 = 2.21e-06  mcrdld_cc_w_40_000_s_10_000 = 3.72e-11  mcrdld_cf_w_40_000_s_10_000 = 1.04e-11
+ mcrdld_ca_w_40_000_s_12_000 = 2.21e-06  mcrdld_cc_w_40_000_s_12_000 = 3.36e-11  mcrdld_cf_w_40_000_s_12_000 = 1.19e-11
+ mcrdld_ca_w_40_000_s_30_000 = 2.21e-06  mcrdld_cc_w_40_000_s_30_000 = 1.82e-11  mcrdld_cf_w_40_000_s_30_000 = 2.15e-11
+ mcrdlp1_ca_w_10_000_s_5_000 = 2.24e-06  mcrdlp1_cc_w_10_000_s_5_000 = 4.08e-11  mcrdlp1_cf_w_10_000_s_5_000 = 6.20e-12
+ mcrdlp1_ca_w_10_000_s_8_000 = 2.24e-06  mcrdlp1_cc_w_10_000_s_8_000 = 3.13e-11  mcrdlp1_cf_w_10_000_s_8_000 = 8.86e-12
+ mcrdlp1_ca_w_10_000_s_10_000 = 2.24e-06  mcrdlp1_cc_w_10_000_s_10_000 = 2.72e-11  mcrdlp1_cf_w_10_000_s_10_000 = 1.05e-11
+ mcrdlp1_ca_w_10_000_s_12_000 = 2.24e-06  mcrdlp1_cc_w_10_000_s_12_000 = 2.40e-11  mcrdlp1_cf_w_10_000_s_12_000 = 1.19e-11
+ mcrdlp1_ca_w_10_000_s_30_000 = 2.24e-06  mcrdlp1_cc_w_10_000_s_30_000 = 1.09e-11  mcrdlp1_cf_w_10_000_s_30_000 = 2.09e-11
+ mcrdlp1_ca_w_40_000_s_5_000 = 2.24e-06  mcrdlp1_cc_w_40_000_s_5_000 = 5.21e-11  mcrdlp1_cf_w_40_000_s_5_000 = 6.30e-12
+ mcrdlp1_ca_w_40_000_s_8_000 = 2.24e-06  mcrdlp1_cc_w_40_000_s_8_000 = 4.16e-11  mcrdlp1_cf_w_40_000_s_8_000 = 8.95e-12
+ mcrdlp1_ca_w_40_000_s_10_000 = 2.24e-06  mcrdlp1_cc_w_40_000_s_10_000 = 3.70e-11  mcrdlp1_cf_w_40_000_s_10_000 = 1.06e-11
+ mcrdlp1_ca_w_40_000_s_12_000 = 2.24e-06  mcrdlp1_cc_w_40_000_s_12_000 = 3.35e-11  mcrdlp1_cf_w_40_000_s_12_000 = 1.21e-11
+ mcrdlp1_ca_w_40_000_s_30_000 = 2.24e-06  mcrdlp1_cc_w_40_000_s_30_000 = 1.81e-11  mcrdlp1_cf_w_40_000_s_30_000 = 2.17e-11
+ mcrdll1_ca_w_10_000_s_5_000 = 2.33e-06  mcrdll1_cc_w_10_000_s_5_000 = 4.05e-11  mcrdll1_cf_w_10_000_s_5_000 = 6.43e-12
+ mcrdll1_ca_w_10_000_s_8_000 = 2.33e-06  mcrdll1_cc_w_10_000_s_8_000 = 3.09e-11  mcrdll1_cf_w_10_000_s_8_000 = 9.16e-12
+ mcrdll1_ca_w_10_000_s_10_000 = 2.33e-06  mcrdll1_cc_w_10_000_s_10_000 = 2.68e-11  mcrdll1_cf_w_10_000_s_10_000 = 1.08e-11
+ mcrdll1_ca_w_10_000_s_12_000 = 2.33e-06  mcrdll1_cc_w_10_000_s_12_000 = 2.37e-11  mcrdll1_cf_w_10_000_s_12_000 = 1.23e-11
+ mcrdll1_ca_w_10_000_s_30_000 = 2.33e-06  mcrdll1_cc_w_10_000_s_30_000 = 1.07e-11  mcrdll1_cf_w_10_000_s_30_000 = 2.13e-11
+ mcrdll1_ca_w_40_000_s_5_000 = 2.33e-06  mcrdll1_cc_w_40_000_s_5_000 = 5.18e-11  mcrdll1_cf_w_40_000_s_5_000 = 6.51e-12
+ mcrdll1_ca_w_40_000_s_8_000 = 2.33e-06  mcrdll1_cc_w_40_000_s_8_000 = 4.13e-11  mcrdll1_cf_w_40_000_s_8_000 = 9.26e-12
+ mcrdll1_ca_w_40_000_s_10_000 = 2.33e-06  mcrdll1_cc_w_40_000_s_10_000 = 3.67e-11  mcrdll1_cf_w_40_000_s_10_000 = 1.09e-11
+ mcrdll1_ca_w_40_000_s_12_000 = 2.33e-06  mcrdll1_cc_w_40_000_s_12_000 = 3.32e-11  mcrdll1_cf_w_40_000_s_12_000 = 1.25e-11
+ mcrdll1_ca_w_40_000_s_30_000 = 2.33e-06  mcrdll1_cc_w_40_000_s_30_000 = 1.78e-11  mcrdll1_cf_w_40_000_s_30_000 = 2.23e-11
+ mcrdlm1_ca_w_10_000_s_5_000 = 2.46e-06  mcrdlm1_cc_w_10_000_s_5_000 = 4.01e-11  mcrdlm1_cf_w_10_000_s_5_000 = 6.75e-12
+ mcrdlm1_ca_w_10_000_s_8_000 = 2.46e-06  mcrdlm1_cc_w_10_000_s_8_000 = 3.05e-11  mcrdlm1_cf_w_10_000_s_8_000 = 9.59e-12
+ mcrdlm1_ca_w_10_000_s_10_000 = 2.46e-06  mcrdlm1_cc_w_10_000_s_10_000 = 2.64e-11  mcrdlm1_cf_w_10_000_s_10_000 = 1.13e-11
+ mcrdlm1_ca_w_10_000_s_12_000 = 2.46e-06  mcrdlm1_cc_w_10_000_s_12_000 = 2.33e-11  mcrdlm1_cf_w_10_000_s_12_000 = 1.29e-11
+ mcrdlm1_ca_w_10_000_s_30_000 = 2.46e-06  mcrdlm1_cc_w_10_000_s_30_000 = 1.04e-11  mcrdlm1_cf_w_10_000_s_30_000 = 2.20e-11
+ mcrdlm1_ca_w_40_000_s_5_000 = 2.46e-06  mcrdlm1_cc_w_40_000_s_5_000 = 5.13e-11  mcrdlm1_cf_w_40_000_s_5_000 = 6.82e-12
+ mcrdlm1_ca_w_40_000_s_8_000 = 2.46e-06  mcrdlm1_cc_w_40_000_s_8_000 = 4.08e-11  mcrdlm1_cf_w_40_000_s_8_000 = 9.67e-12
+ mcrdlm1_ca_w_40_000_s_10_000 = 2.46e-06  mcrdlm1_cc_w_40_000_s_10_000 = 3.62e-11  mcrdlm1_cf_w_40_000_s_10_000 = 1.14e-11
+ mcrdlm1_ca_w_40_000_s_12_000 = 2.46e-06  mcrdlm1_cc_w_40_000_s_12_000 = 3.27e-11  mcrdlm1_cf_w_40_000_s_12_000 = 1.30e-11
+ mcrdlm1_ca_w_40_000_s_30_000 = 2.46e-06  mcrdlm1_cc_w_40_000_s_30_000 = 1.75e-11  mcrdlm1_cf_w_40_000_s_30_000 = 2.29e-11
+ mcrdlm2_ca_w_10_000_s_5_000 = 2.60e-06  mcrdlm2_cc_w_10_000_s_5_000 = 3.96e-11  mcrdlm2_cf_w_10_000_s_5_000 = 7.09e-12
+ mcrdlm2_ca_w_10_000_s_8_000 = 2.60e-06  mcrdlm2_cc_w_10_000_s_8_000 = 3.00e-11  mcrdlm2_cf_w_10_000_s_8_000 = 1.01e-11
+ mcrdlm2_ca_w_10_000_s_10_000 = 2.60e-06  mcrdlm2_cc_w_10_000_s_10_000 = 2.59e-11  mcrdlm2_cf_w_10_000_s_10_000 = 1.18e-11
+ mcrdlm2_ca_w_10_000_s_12_000 = 2.60e-06  mcrdlm2_cc_w_10_000_s_12_000 = 2.28e-11  mcrdlm2_cf_w_10_000_s_12_000 = 1.34e-11
+ mcrdlm2_ca_w_10_000_s_30_000 = 2.60e-06  mcrdlm2_cc_w_10_000_s_30_000 = 1.00e-11  mcrdlm2_cf_w_10_000_s_30_000 = 2.26e-11
+ mcrdlm2_ca_w_40_000_s_5_000 = 2.60e-06  mcrdlm2_cc_w_40_000_s_5_000 = 5.08e-11  mcrdlm2_cf_w_40_000_s_5_000 = 7.16e-12
+ mcrdlm2_ca_w_40_000_s_8_000 = 2.60e-06  mcrdlm2_cc_w_40_000_s_8_000 = 4.02e-11  mcrdlm2_cf_w_40_000_s_8_000 = 1.01e-11
+ mcrdlm2_ca_w_40_000_s_10_000 = 2.60e-06  mcrdlm2_cc_w_40_000_s_10_000 = 3.58e-11  mcrdlm2_cf_w_40_000_s_10_000 = 1.19e-11
+ mcrdlm2_ca_w_40_000_s_12_000 = 2.60e-06  mcrdlm2_cc_w_40_000_s_12_000 = 3.23e-11  mcrdlm2_cf_w_40_000_s_12_000 = 1.36e-11
+ mcrdlm2_ca_w_40_000_s_30_000 = 2.60e-06  mcrdlm2_cc_w_40_000_s_30_000 = 1.72e-11  mcrdlm2_cf_w_40_000_s_30_000 = 2.37e-11
+ mcrdlm3_ca_w_10_000_s_5_000 = 2.90e-06  mcrdlm3_cc_w_10_000_s_5_000 = 3.87e-11  mcrdlm3_cf_w_10_000_s_5_000 = 7.76e-12
+ mcrdlm3_ca_w_10_000_s_8_000 = 2.90e-06  mcrdlm3_cc_w_10_000_s_8_000 = 2.91e-11  mcrdlm3_cf_w_10_000_s_8_000 = 1.09e-11
+ mcrdlm3_ca_w_10_000_s_10_000 = 2.90e-06  mcrdlm3_cc_w_10_000_s_10_000 = 2.51e-11  mcrdlm3_cf_w_10_000_s_10_000 = 1.28e-11
+ mcrdlm3_ca_w_10_000_s_12_000 = 2.90e-06  mcrdlm3_cc_w_10_000_s_12_000 = 2.20e-11  mcrdlm3_cf_w_10_000_s_12_000 = 1.45e-11
+ mcrdlm3_ca_w_10_000_s_30_000 = 2.90e-06  mcrdlm3_cc_w_10_000_s_30_000 = 9.43e-12  mcrdlm3_cf_w_10_000_s_30_000 = 2.39e-11
+ mcrdlm3_ca_w_40_000_s_5_000 = 2.90e-06  mcrdlm3_cc_w_40_000_s_5_000 = 4.99e-11  mcrdlm3_cf_w_40_000_s_5_000 = 7.73e-12
+ mcrdlm3_ca_w_40_000_s_8_000 = 2.90e-06  mcrdlm3_cc_w_40_000_s_8_000 = 3.94e-11  mcrdlm3_cf_w_40_000_s_8_000 = 1.09e-11
+ mcrdlm3_ca_w_40_000_s_10_000 = 2.90e-06  mcrdlm3_cc_w_40_000_s_10_000 = 3.49e-11  mcrdlm3_cf_w_40_000_s_10_000 = 1.28e-11
+ mcrdlm3_ca_w_40_000_s_12_000 = 2.90e-06  mcrdlm3_cc_w_40_000_s_12_000 = 3.14e-11  mcrdlm3_cf_w_40_000_s_12_000 = 1.46e-11
+ mcrdlm3_ca_w_40_000_s_30_000 = 2.90e-06  mcrdlm3_cc_w_40_000_s_30_000 = 1.65e-11  mcrdlm3_cf_w_40_000_s_30_000 = 2.49e-11
+ mcrdlm4_ca_w_10_000_s_5_000 = 3.28e-06  mcrdlm4_cc_w_10_000_s_5_000 = 3.78e-11  mcrdlm4_cf_w_10_000_s_5_000 = 8.63e-12
+ mcrdlm4_ca_w_10_000_s_8_000 = 3.28e-06  mcrdlm4_cc_w_10_000_s_8_000 = 2.82e-11  mcrdlm4_cf_w_10_000_s_8_000 = 1.21e-11
+ mcrdlm4_ca_w_10_000_s_10_000 = 3.28e-06  mcrdlm4_cc_w_10_000_s_10_000 = 2.42e-11  mcrdlm4_cf_w_10_000_s_10_000 = 1.41e-11
+ mcrdlm4_ca_w_10_000_s_12_000 = 3.28e-06  mcrdlm4_cc_w_10_000_s_12_000 = 2.11e-11  mcrdlm4_cf_w_10_000_s_12_000 = 1.59e-11
+ mcrdlm4_ca_w_10_000_s_30_000 = 3.28e-06  mcrdlm4_cc_w_10_000_s_30_000 = 8.80e-12  mcrdlm4_cf_w_10_000_s_30_000 = 2.54e-11
+ mcrdlm4_ca_w_40_000_s_5_000 = 3.28e-06  mcrdlm4_cc_w_40_000_s_5_000 = 4.89e-11  mcrdlm4_cf_w_40_000_s_5_000 = 8.55e-12
+ mcrdlm4_ca_w_40_000_s_8_000 = 3.28e-06  mcrdlm4_cc_w_40_000_s_8_000 = 3.85e-11  mcrdlm4_cf_w_40_000_s_8_000 = 1.20e-11
+ mcrdlm4_ca_w_40_000_s_10_000 = 3.28e-06  mcrdlm4_cc_w_40_000_s_10_000 = 3.39e-11  mcrdlm4_cf_w_40_000_s_10_000 = 1.41e-11
+ mcrdlm4_ca_w_40_000_s_12_000 = 3.28e-06  mcrdlm4_cc_w_40_000_s_12_000 = 3.05e-11  mcrdlm4_cf_w_40_000_s_12_000 = 1.59e-11
+ mcrdlm4_ca_w_40_000_s_30_000 = 3.28e-06  mcrdlm4_cc_w_40_000_s_30_000 = 1.59e-11  mcrdlm4_cf_w_40_000_s_30_000 = 2.64e-11
+ mcrdlm5_ca_w_10_000_s_5_000 = 4.28e-06  mcrdlm5_cc_w_10_000_s_5_000 = 3.57e-11  mcrdlm5_cf_w_10_000_s_5_000 = 1.09e-11
+ mcrdlm5_ca_w_10_000_s_8_000 = 4.28e-06  mcrdlm5_cc_w_10_000_s_8_000 = 2.62e-11  mcrdlm5_cf_w_10_000_s_8_000 = 1.49e-11
+ mcrdlm5_ca_w_10_000_s_10_000 = 4.28e-06  mcrdlm5_cc_w_10_000_s_10_000 = 2.22e-11  mcrdlm5_cf_w_10_000_s_10_000 = 1.72e-11
+ mcrdlm5_ca_w_10_000_s_12_000 = 4.28e-06  mcrdlm5_cc_w_10_000_s_12_000 = 1.92e-11  mcrdlm5_cf_w_10_000_s_12_000 = 1.91e-11
+ mcrdlm5_ca_w_10_000_s_30_000 = 4.28e-06  mcrdlm5_cc_w_10_000_s_30_000 = 7.63e-12  mcrdlm5_cf_w_10_000_s_30_000 = 2.86e-11
+ mcrdlm5_ca_w_40_000_s_5_000 = 4.28e-06  mcrdlm5_cc_w_40_000_s_5_000 = 4.67e-11  mcrdlm5_cf_w_40_000_s_5_000 = 1.08e-11
+ mcrdlm5_ca_w_40_000_s_8_000 = 4.28e-06  mcrdlm5_cc_w_40_000_s_8_000 = 3.64e-11  mcrdlm5_cf_w_40_000_s_8_000 = 1.48e-11
+ mcrdlm5_ca_w_40_000_s_10_000 = 4.28e-06  mcrdlm5_cc_w_40_000_s_10_000 = 3.20e-11  mcrdlm5_cf_w_40_000_s_10_000 = 1.72e-11
+ mcrdlm5_ca_w_40_000_s_12_000 = 4.28e-06  mcrdlm5_cc_w_40_000_s_12_000 = 2.87e-11  mcrdlm5_cf_w_40_000_s_12_000 = 1.92e-11
+ mcrdlm5_ca_w_40_000_s_30_000 = 4.28e-06  mcrdlm5_cc_w_40_000_s_30_000 = 1.46e-11  mcrdlm5_cf_w_40_000_s_30_000 = 3.01e-11
+ mcl1p1f_ca_w_0_150_s_0_210 = 1.45e-04  mcl1p1f_cc_w_0_150_s_0_210 = 5.70e-11  mcl1p1f_cf_w_0_150_s_0_210 = 1.54e-11
+ mcl1p1f_ca_w_0_150_s_0_263 = 1.45e-04  mcl1p1f_cc_w_0_150_s_0_263 = 4.57e-11  mcl1p1f_cf_w_0_150_s_0_263 = 1.85e-11
+ mcl1p1f_ca_w_0_150_s_0_315 = 1.45e-04  mcl1p1f_cc_w_0_150_s_0_315 = 3.74e-11  mcl1p1f_cf_w_0_150_s_0_315 = 2.13e-11
+ mcl1p1f_ca_w_0_150_s_0_420 = 1.45e-04  mcl1p1f_cc_w_0_150_s_0_420 = 2.65e-11  mcl1p1f_cf_w_0_150_s_0_420 = 2.64e-11
+ mcl1p1f_ca_w_0_150_s_0_525 = 1.45e-04  mcl1p1f_cc_w_0_150_s_0_525 = 1.92e-11  mcl1p1f_cf_w_0_150_s_0_525 = 3.05e-11
+ mcl1p1f_ca_w_0_150_s_0_630 = 1.45e-04  mcl1p1f_cc_w_0_150_s_0_630 = 1.42e-11  mcl1p1f_cf_w_0_150_s_0_630 = 3.39e-11
+ mcl1p1f_ca_w_0_150_s_0_840 = 1.45e-04  mcl1p1f_cc_w_0_150_s_0_840 = 7.96e-12  mcl1p1f_cf_w_0_150_s_0_840 = 3.88e-11
+ mcl1p1f_ca_w_0_150_s_1_260 = 1.45e-04  mcl1p1f_cc_w_0_150_s_1_260 = 2.59e-12  mcl1p1f_cf_w_0_150_s_1_260 = 4.37e-11
+ mcl1p1f_ca_w_0_150_s_2_310 = 1.45e-04  mcl1p1f_cc_w_0_150_s_2_310 = 1.95e-13  mcl1p1f_cf_w_0_150_s_2_310 = 4.59e-11
+ mcl1p1f_ca_w_0_150_s_5_250 = 1.45e-04  mcl1p1f_cc_w_0_150_s_5_250 = 3.23e-27  mcl1p1f_cf_w_0_150_s_5_250 = 4.62e-11
+ mcl1p1f_ca_w_1_200_s_0_210 = 1.45e-04  mcl1p1f_cc_w_1_200_s_0_210 = 6.11e-11  mcl1p1f_cf_w_1_200_s_0_210 = 1.54e-11
+ mcl1p1f_ca_w_1_200_s_0_263 = 1.45e-04  mcl1p1f_cc_w_1_200_s_0_263 = 4.88e-11  mcl1p1f_cf_w_1_200_s_0_263 = 1.85e-11
+ mcl1p1f_ca_w_1_200_s_0_315 = 1.45e-04  mcl1p1f_cc_w_1_200_s_0_315 = 4.02e-11  mcl1p1f_cf_w_1_200_s_0_315 = 2.13e-11
+ mcl1p1f_ca_w_1_200_s_0_420 = 1.45e-04  mcl1p1f_cc_w_1_200_s_0_420 = 2.85e-11  mcl1p1f_cf_w_1_200_s_0_420 = 2.65e-11
+ mcl1p1f_ca_w_1_200_s_0_525 = 1.45e-04  mcl1p1f_cc_w_1_200_s_0_525 = 2.09e-11  mcl1p1f_cf_w_1_200_s_0_525 = 3.09e-11
+ mcl1p1f_ca_w_1_200_s_0_630 = 1.45e-04  mcl1p1f_cc_w_1_200_s_0_630 = 1.54e-11  mcl1p1f_cf_w_1_200_s_0_630 = 3.45e-11
+ mcl1p1f_ca_w_1_200_s_0_840 = 1.45e-04  mcl1p1f_cc_w_1_200_s_0_840 = 8.75e-12  mcl1p1f_cf_w_1_200_s_0_840 = 3.97e-11
+ mcl1p1f_ca_w_1_200_s_1_260 = 1.45e-04  mcl1p1f_cc_w_1_200_s_1_260 = 2.90e-12  mcl1p1f_cf_w_1_200_s_1_260 = 4.49e-11
+ mcl1p1f_ca_w_1_200_s_2_310 = 1.45e-04  mcl1p1f_cc_w_1_200_s_2_310 = 2.00e-13  mcl1p1f_cf_w_1_200_s_2_310 = 4.74e-11
+ mcl1p1f_ca_w_1_200_s_5_250 = 1.45e-04  mcl1p1f_cc_w_1_200_s_5_250 = 0.00e+00  mcl1p1f_cf_w_1_200_s_5_250 = 4.76e-11
+ mcm1p1f_ca_w_0_150_s_0_210 = 1.13e-04  mcm1p1f_cc_w_0_150_s_0_210 = 6.11e-11  mcm1p1f_cf_w_0_150_s_0_210 = 1.22e-11
+ mcm1p1f_ca_w_0_150_s_0_263 = 1.13e-04  mcm1p1f_cc_w_0_150_s_0_263 = 5.00e-11  mcm1p1f_cf_w_0_150_s_0_263 = 1.46e-11
+ mcm1p1f_ca_w_0_150_s_0_315 = 1.13e-04  mcm1p1f_cc_w_0_150_s_0_315 = 4.20e-11  mcm1p1f_cf_w_0_150_s_0_315 = 1.69e-11
+ mcm1p1f_ca_w_0_150_s_0_420 = 1.13e-04  mcm1p1f_cc_w_0_150_s_0_420 = 3.13e-11  mcm1p1f_cf_w_0_150_s_0_420 = 2.12e-11
+ mcm1p1f_ca_w_0_150_s_0_525 = 1.13e-04  mcm1p1f_cc_w_0_150_s_0_525 = 2.41e-11  mcm1p1f_cf_w_0_150_s_0_525 = 2.49e-11
+ mcm1p1f_ca_w_0_150_s_0_630 = 1.13e-04  mcm1p1f_cc_w_0_150_s_0_630 = 1.89e-11  mcm1p1f_cf_w_0_150_s_0_630 = 2.80e-11
+ mcm1p1f_ca_w_0_150_s_0_840 = 1.13e-04  mcm1p1f_cc_w_0_150_s_0_840 = 1.21e-11  mcm1p1f_cf_w_0_150_s_0_840 = 3.28e-11
+ mcm1p1f_ca_w_0_150_s_1_260 = 1.13e-04  mcm1p1f_cc_w_0_150_s_1_260 = 5.24e-12  mcm1p1f_cf_w_0_150_s_1_260 = 3.85e-11
+ mcm1p1f_ca_w_0_150_s_2_310 = 1.13e-04  mcm1p1f_cc_w_0_150_s_2_310 = 7.85e-13  mcm1p1f_cf_w_0_150_s_2_310 = 4.26e-11
+ mcm1p1f_ca_w_0_150_s_5_250 = 1.13e-04  mcm1p1f_cc_w_0_150_s_5_250 = 2.00e-14  mcm1p1f_cf_w_0_150_s_5_250 = 4.34e-11
+ mcm1p1f_ca_w_1_200_s_0_210 = 1.13e-04  mcm1p1f_cc_w_1_200_s_0_210 = 6.86e-11  mcm1p1f_cf_w_1_200_s_0_210 = 1.21e-11
+ mcm1p1f_ca_w_1_200_s_0_263 = 1.13e-04  mcm1p1f_cc_w_1_200_s_0_263 = 5.64e-11  mcm1p1f_cf_w_1_200_s_0_263 = 1.47e-11
+ mcm1p1f_ca_w_1_200_s_0_315 = 1.13e-04  mcm1p1f_cc_w_1_200_s_0_315 = 4.77e-11  mcm1p1f_cf_w_1_200_s_0_315 = 1.70e-11
+ mcm1p1f_ca_w_1_200_s_0_420 = 1.13e-04  mcm1p1f_cc_w_1_200_s_0_420 = 3.58e-11  mcm1p1f_cf_w_1_200_s_0_420 = 2.13e-11
+ mcm1p1f_ca_w_1_200_s_0_525 = 1.13e-04  mcm1p1f_cc_w_1_200_s_0_525 = 2.78e-11  mcm1p1f_cf_w_1_200_s_0_525 = 2.52e-11
+ mcm1p1f_ca_w_1_200_s_0_630 = 1.13e-04  mcm1p1f_cc_w_1_200_s_0_630 = 2.20e-11  mcm1p1f_cf_w_1_200_s_0_630 = 2.85e-11
+ mcm1p1f_ca_w_1_200_s_0_840 = 1.13e-04  mcm1p1f_cc_w_1_200_s_0_840 = 1.43e-11  mcm1p1f_cf_w_1_200_s_0_840 = 3.37e-11
+ mcm1p1f_ca_w_1_200_s_1_260 = 1.13e-04  mcm1p1f_cc_w_1_200_s_1_260 = 6.41e-12  mcm1p1f_cf_w_1_200_s_1_260 = 4.01e-11
+ mcm1p1f_ca_w_1_200_s_2_310 = 1.13e-04  mcm1p1f_cc_w_1_200_s_2_310 = 1.03e-12  mcm1p1f_cf_w_1_200_s_2_310 = 4.52e-11
+ mcm1p1f_ca_w_1_200_s_5_250 = 1.13e-04  mcm1p1f_cc_w_1_200_s_5_250 = 5.00e-14  mcm1p1f_cf_w_1_200_s_5_250 = 4.62e-11
+ mcm2p1f_ca_w_0_150_s_0_210 = 9.94e-05  mcm2p1f_cc_w_0_150_s_0_210 = 6.30e-11  mcm2p1f_cf_w_0_150_s_0_210 = 1.08e-11
+ mcm2p1f_ca_w_0_150_s_0_263 = 9.94e-05  mcm2p1f_cc_w_0_150_s_0_263 = 5.20e-11  mcm2p1f_cf_w_0_150_s_0_263 = 1.29e-11
+ mcm2p1f_ca_w_0_150_s_0_315 = 9.94e-05  mcm2p1f_cc_w_0_150_s_0_315 = 4.44e-11  mcm2p1f_cf_w_0_150_s_0_315 = 1.50e-11
+ mcm2p1f_ca_w_0_150_s_0_420 = 9.94e-05  mcm2p1f_cc_w_0_150_s_0_420 = 3.38e-11  mcm2p1f_cf_w_0_150_s_0_420 = 1.88e-11
+ mcm2p1f_ca_w_0_150_s_0_525 = 9.94e-05  mcm2p1f_cc_w_0_150_s_0_525 = 2.68e-11  mcm2p1f_cf_w_0_150_s_0_525 = 2.21e-11
+ mcm2p1f_ca_w_0_150_s_0_630 = 9.94e-05  mcm2p1f_cc_w_0_150_s_0_630 = 2.18e-11  mcm2p1f_cf_w_0_150_s_0_630 = 2.50e-11
+ mcm2p1f_ca_w_0_150_s_0_840 = 9.94e-05  mcm2p1f_cc_w_0_150_s_0_840 = 1.48e-11  mcm2p1f_cf_w_0_150_s_0_840 = 2.97e-11
+ mcm2p1f_ca_w_0_150_s_1_260 = 9.94e-05  mcm2p1f_cc_w_0_150_s_1_260 = 7.41e-12  mcm2p1f_cf_w_0_150_s_1_260 = 3.56e-11
+ mcm2p1f_ca_w_0_150_s_2_310 = 9.94e-05  mcm2p1f_cc_w_0_150_s_2_310 = 1.71e-12  mcm2p1f_cf_w_0_150_s_2_310 = 4.08e-11
+ mcm2p1f_ca_w_0_150_s_5_250 = 9.94e-05  mcm2p1f_cc_w_0_150_s_5_250 = 8.00e-14  mcm2p1f_cf_w_0_150_s_5_250 = 4.24e-11
+ mcm2p1f_ca_w_1_200_s_0_210 = 9.94e-05  mcm2p1f_cc_w_1_200_s_0_210 = 7.39e-11  mcm2p1f_cf_w_1_200_s_0_210 = 1.07e-11
+ mcm2p1f_ca_w_1_200_s_0_263 = 9.94e-05  mcm2p1f_cc_w_1_200_s_0_263 = 6.16e-11  mcm2p1f_cf_w_1_200_s_0_263 = 1.30e-11
+ mcm2p1f_ca_w_1_200_s_0_315 = 9.94e-05  mcm2p1f_cc_w_1_200_s_0_315 = 5.30e-11  mcm2p1f_cf_w_1_200_s_0_315 = 1.50e-11
+ mcm2p1f_ca_w_1_200_s_0_420 = 9.94e-05  mcm2p1f_cc_w_1_200_s_0_420 = 4.11e-11  mcm2p1f_cf_w_1_200_s_0_420 = 1.89e-11
+ mcm2p1f_ca_w_1_200_s_0_525 = 9.94e-05  mcm2p1f_cc_w_1_200_s_0_525 = 3.30e-11  mcm2p1f_cf_w_1_200_s_0_525 = 2.24e-11
+ mcm2p1f_ca_w_1_200_s_0_630 = 9.94e-05  mcm2p1f_cc_w_1_200_s_0_630 = 2.72e-11  mcm2p1f_cf_w_1_200_s_0_630 = 2.54e-11
+ mcm2p1f_ca_w_1_200_s_0_840 = 9.94e-05  mcm2p1f_cc_w_1_200_s_0_840 = 1.91e-11  mcm2p1f_cf_w_1_200_s_0_840 = 3.05e-11
+ mcm2p1f_ca_w_1_200_s_1_260 = 9.94e-05  mcm2p1f_cc_w_1_200_s_1_260 = 1.02e-11  mcm2p1f_cf_w_1_200_s_1_260 = 3.73e-11
+ mcm2p1f_ca_w_1_200_s_2_310 = 9.94e-05  mcm2p1f_cc_w_1_200_s_2_310 = 2.59e-12  mcm2p1f_cf_w_1_200_s_2_310 = 4.41e-11
+ mcm2p1f_ca_w_1_200_s_5_250 = 9.94e-05  mcm2p1f_cc_w_1_200_s_5_250 = 1.15e-13  mcm2p1f_cf_w_1_200_s_5_250 = 4.65e-11
+ mcm3p1f_ca_w_0_150_s_0_210 = 9.31e-05  mcm3p1f_cc_w_0_150_s_0_210 = 6.39e-11  mcm3p1f_cf_w_0_150_s_0_210 = 1.01e-11
+ mcm3p1f_ca_w_0_150_s_0_263 = 9.31e-05  mcm3p1f_cc_w_0_150_s_0_263 = 5.30e-11  mcm3p1f_cf_w_0_150_s_0_263 = 1.21e-11
+ mcm3p1f_ca_w_0_150_s_0_315 = 9.31e-05  mcm3p1f_cc_w_0_150_s_0_315 = 4.56e-11  mcm3p1f_cf_w_0_150_s_0_315 = 1.40e-11
+ mcm3p1f_ca_w_0_150_s_0_420 = 9.31e-05  mcm3p1f_cc_w_0_150_s_0_420 = 3.51e-11  mcm3p1f_cf_w_0_150_s_0_420 = 1.77e-11
+ mcm3p1f_ca_w_0_150_s_0_525 = 9.31e-05  mcm3p1f_cc_w_0_150_s_0_525 = 2.83e-11  mcm3p1f_cf_w_0_150_s_0_525 = 2.08e-11
+ mcm3p1f_ca_w_0_150_s_0_630 = 9.31e-05  mcm3p1f_cc_w_0_150_s_0_630 = 2.33e-11  mcm3p1f_cf_w_0_150_s_0_630 = 2.35e-11
+ mcm3p1f_ca_w_0_150_s_0_840 = 9.31e-05  mcm3p1f_cc_w_0_150_s_0_840 = 1.64e-11  mcm3p1f_cf_w_0_150_s_0_840 = 2.81e-11
+ mcm3p1f_ca_w_0_150_s_1_260 = 9.31e-05  mcm3p1f_cc_w_0_150_s_1_260 = 8.77e-12  mcm3p1f_cf_w_0_150_s_1_260 = 3.41e-11
+ mcm3p1f_ca_w_0_150_s_2_310 = 9.31e-05  mcm3p1f_cc_w_0_150_s_2_310 = 2.52e-12  mcm3p1f_cf_w_0_150_s_2_310 = 3.97e-11
+ mcm3p1f_ca_w_0_150_s_5_250 = 9.31e-05  mcm3p1f_cc_w_0_150_s_5_250 = 1.85e-13  mcm3p1f_cf_w_0_150_s_5_250 = 4.20e-11
+ mcm3p1f_ca_w_1_200_s_0_210 = 9.31e-05  mcm3p1f_cc_w_1_200_s_0_210 = 7.69e-11  mcm3p1f_cf_w_1_200_s_0_210 = 1.00e-11
+ mcm3p1f_ca_w_1_200_s_0_263 = 9.31e-05  mcm3p1f_cc_w_1_200_s_0_263 = 6.48e-11  mcm3p1f_cf_w_1_200_s_0_263 = 1.21e-11
+ mcm3p1f_ca_w_1_200_s_0_315 = 9.31e-05  mcm3p1f_cc_w_1_200_s_0_315 = 5.62e-11  mcm3p1f_cf_w_1_200_s_0_315 = 1.41e-11
+ mcm3p1f_ca_w_1_200_s_0_420 = 9.31e-05  mcm3p1f_cc_w_1_200_s_0_420 = 4.44e-11  mcm3p1f_cf_w_1_200_s_0_420 = 1.77e-11
+ mcm3p1f_ca_w_1_200_s_0_525 = 9.31e-05  mcm3p1f_cc_w_1_200_s_0_525 = 3.64e-11  mcm3p1f_cf_w_1_200_s_0_525 = 2.10e-11
+ mcm3p1f_ca_w_1_200_s_0_630 = 9.31e-05  mcm3p1f_cc_w_1_200_s_0_630 = 3.04e-11  mcm3p1f_cf_w_1_200_s_0_630 = 2.39e-11
+ mcm3p1f_ca_w_1_200_s_0_840 = 9.31e-05  mcm3p1f_cc_w_1_200_s_0_840 = 2.23e-11  mcm3p1f_cf_w_1_200_s_0_840 = 2.88e-11
+ mcm3p1f_ca_w_1_200_s_1_260 = 9.31e-05  mcm3p1f_cc_w_1_200_s_1_260 = 1.31e-11  mcm3p1f_cf_w_1_200_s_1_260 = 3.56e-11
+ mcm3p1f_ca_w_1_200_s_2_310 = 9.31e-05  mcm3p1f_cc_w_1_200_s_2_310 = 4.17e-12  mcm3p1f_cf_w_1_200_s_2_310 = 4.33e-11
+ mcm3p1f_ca_w_1_200_s_5_250 = 9.31e-05  mcm3p1f_cc_w_1_200_s_5_250 = 2.95e-13  mcm3p1f_cf_w_1_200_s_5_250 = 4.71e-11
+ mcm4p1f_ca_w_0_150_s_0_210 = 8.89e-05  mcm4p1f_cc_w_0_150_s_0_210 = 6.45e-11  mcm4p1f_cf_w_0_150_s_0_210 = 9.64e-12
+ mcm4p1f_ca_w_0_150_s_0_263 = 8.89e-05  mcm4p1f_cc_w_0_150_s_0_263 = 5.37e-11  mcm4p1f_cf_w_0_150_s_0_263 = 1.15e-11
+ mcm4p1f_ca_w_0_150_s_0_315 = 8.89e-05  mcm4p1f_cc_w_0_150_s_0_315 = 4.64e-11  mcm4p1f_cf_w_0_150_s_0_315 = 1.33e-11
+ mcm4p1f_ca_w_0_150_s_0_420 = 8.89e-05  mcm4p1f_cc_w_0_150_s_0_420 = 3.60e-11  mcm4p1f_cf_w_0_150_s_0_420 = 1.69e-11
+ mcm4p1f_ca_w_0_150_s_0_525 = 8.89e-05  mcm4p1f_cc_w_0_150_s_0_525 = 2.93e-11  mcm4p1f_cf_w_0_150_s_0_525 = 1.98e-11
+ mcm4p1f_ca_w_0_150_s_0_630 = 8.89e-05  mcm4p1f_cc_w_0_150_s_0_630 = 2.44e-11  mcm4p1f_cf_w_0_150_s_0_630 = 2.25e-11
+ mcm4p1f_ca_w_0_150_s_0_840 = 8.89e-05  mcm4p1f_cc_w_0_150_s_0_840 = 1.76e-11  mcm4p1f_cf_w_0_150_s_0_840 = 2.69e-11
+ mcm4p1f_ca_w_0_150_s_1_260 = 8.89e-05  mcm4p1f_cc_w_0_150_s_1_260 = 9.77e-12  mcm4p1f_cf_w_0_150_s_1_260 = 3.31e-11
+ mcm4p1f_ca_w_0_150_s_2_310 = 8.89e-05  mcm4p1f_cc_w_0_150_s_2_310 = 3.26e-12  mcm4p1f_cf_w_0_150_s_2_310 = 3.88e-11
+ mcm4p1f_ca_w_0_150_s_5_250 = 8.89e-05  mcm4p1f_cc_w_0_150_s_5_250 = 3.70e-13  mcm4p1f_cf_w_0_150_s_5_250 = 4.17e-11
+ mcm4p1f_ca_w_1_200_s_0_210 = 8.89e-05  mcm4p1f_cc_w_1_200_s_0_210 = 7.92e-11  mcm4p1f_cf_w_1_200_s_0_210 = 9.57e-12
+ mcm4p1f_ca_w_1_200_s_0_263 = 8.89e-05  mcm4p1f_cc_w_1_200_s_0_263 = 6.72e-11  mcm4p1f_cf_w_1_200_s_0_263 = 1.16e-11
+ mcm4p1f_ca_w_1_200_s_0_315 = 8.89e-05  mcm4p1f_cc_w_1_200_s_0_315 = 5.87e-11  mcm4p1f_cf_w_1_200_s_0_315 = 1.34e-11
+ mcm4p1f_ca_w_1_200_s_0_420 = 8.89e-05  mcm4p1f_cc_w_1_200_s_0_420 = 4.69e-11  mcm4p1f_cf_w_1_200_s_0_420 = 1.69e-11
+ mcm4p1f_ca_w_1_200_s_0_525 = 8.89e-05  mcm4p1f_cc_w_1_200_s_0_525 = 3.89e-11  mcm4p1f_cf_w_1_200_s_0_525 = 2.00e-11
+ mcm4p1f_ca_w_1_200_s_0_630 = 8.89e-05  mcm4p1f_cc_w_1_200_s_0_630 = 3.30e-11  mcm4p1f_cf_w_1_200_s_0_630 = 2.29e-11
+ mcm4p1f_ca_w_1_200_s_0_840 = 8.89e-05  mcm4p1f_cc_w_1_200_s_0_840 = 2.49e-11  mcm4p1f_cf_w_1_200_s_0_840 = 2.76e-11
+ mcm4p1f_ca_w_1_200_s_1_260 = 8.89e-05  mcm4p1f_cc_w_1_200_s_1_260 = 1.54e-11  mcm4p1f_cf_w_1_200_s_1_260 = 3.44e-11
+ mcm4p1f_ca_w_1_200_s_2_310 = 8.89e-05  mcm4p1f_cc_w_1_200_s_2_310 = 5.87e-12  mcm4p1f_cf_w_1_200_s_2_310 = 4.27e-11
+ mcm4p1f_ca_w_1_200_s_5_250 = 8.89e-05  mcm4p1f_cc_w_1_200_s_5_250 = 6.90e-13  mcm4p1f_cf_w_1_200_s_5_250 = 4.76e-11
+ mcm5p1f_ca_w_0_150_s_0_210 = 8.66e-05  mcm5p1f_cc_w_0_150_s_0_210 = 6.48e-11  mcm5p1f_cf_w_0_150_s_0_210 = 9.39e-12
+ mcm5p1f_ca_w_0_150_s_0_263 = 8.66e-05  mcm5p1f_cc_w_0_150_s_0_263 = 5.41e-11  mcm5p1f_cf_w_0_150_s_0_263 = 1.12e-11
+ mcm5p1f_ca_w_0_150_s_0_315 = 8.66e-05  mcm5p1f_cc_w_0_150_s_0_315 = 4.68e-11  mcm5p1f_cf_w_0_150_s_0_315 = 1.30e-11
+ mcm5p1f_ca_w_0_150_s_0_420 = 8.66e-05  mcm5p1f_cc_w_0_150_s_0_420 = 3.64e-11  mcm5p1f_cf_w_0_150_s_0_420 = 1.64e-11
+ mcm5p1f_ca_w_0_150_s_0_525 = 8.66e-05  mcm5p1f_cc_w_0_150_s_0_525 = 2.98e-11  mcm5p1f_cf_w_0_150_s_0_525 = 1.93e-11
+ mcm5p1f_ca_w_0_150_s_0_630 = 8.66e-05  mcm5p1f_cc_w_0_150_s_0_630 = 2.50e-11  mcm5p1f_cf_w_0_150_s_0_630 = 2.19e-11
+ mcm5p1f_ca_w_0_150_s_0_840 = 8.66e-05  mcm5p1f_cc_w_0_150_s_0_840 = 1.82e-11  mcm5p1f_cf_w_0_150_s_0_840 = 2.63e-11
+ mcm5p1f_ca_w_0_150_s_1_260 = 8.66e-05  mcm5p1f_cc_w_0_150_s_1_260 = 1.04e-11  mcm5p1f_cf_w_0_150_s_1_260 = 3.25e-11
+ mcm5p1f_ca_w_0_150_s_2_310 = 8.66e-05  mcm5p1f_cc_w_0_150_s_2_310 = 3.76e-12  mcm5p1f_cf_w_0_150_s_2_310 = 3.83e-11
+ mcm5p1f_ca_w_0_150_s_5_250 = 8.66e-05  mcm5p1f_cc_w_0_150_s_5_250 = 5.27e-13  mcm5p1f_cf_w_0_150_s_5_250 = 4.15e-11
+ mcm5p1f_ca_w_1_200_s_0_210 = 8.66e-05  mcm5p1f_cc_w_1_200_s_0_210 = 8.04e-11  mcm5p1f_cf_w_1_200_s_0_210 = 9.32e-12
+ mcm5p1f_ca_w_1_200_s_0_263 = 8.66e-05  mcm5p1f_cc_w_1_200_s_0_263 = 6.85e-11  mcm5p1f_cf_w_1_200_s_0_263 = 1.12e-11
+ mcm5p1f_ca_w_1_200_s_0_315 = 8.66e-05  mcm5p1f_cc_w_1_200_s_0_315 = 6.00e-11  mcm5p1f_cf_w_1_200_s_0_315 = 1.31e-11
+ mcm5p1f_ca_w_1_200_s_0_420 = 8.66e-05  mcm5p1f_cc_w_1_200_s_0_420 = 4.83e-11  mcm5p1f_cf_w_1_200_s_0_420 = 1.65e-11
+ mcm5p1f_ca_w_1_200_s_0_525 = 8.66e-05  mcm5p1f_cc_w_1_200_s_0_525 = 4.04e-11  mcm5p1f_cf_w_1_200_s_0_525 = 1.95e-11
+ mcm5p1f_ca_w_1_200_s_0_630 = 8.66e-05  mcm5p1f_cc_w_1_200_s_0_630 = 3.45e-11  mcm5p1f_cf_w_1_200_s_0_630 = 2.23e-11
+ mcm5p1f_ca_w_1_200_s_0_840 = 8.66e-05  mcm5p1f_cc_w_1_200_s_0_840 = 2.65e-11  mcm5p1f_cf_w_1_200_s_0_840 = 2.70e-11
+ mcm5p1f_ca_w_1_200_s_1_260 = 8.66e-05  mcm5p1f_cc_w_1_200_s_1_260 = 1.69e-11  mcm5p1f_cf_w_1_200_s_1_260 = 3.37e-11
+ mcm5p1f_ca_w_1_200_s_2_310 = 8.66e-05  mcm5p1f_cc_w_1_200_s_2_310 = 7.02e-12  mcm5p1f_cf_w_1_200_s_2_310 = 4.22e-11
+ mcm5p1f_ca_w_1_200_s_5_250 = 8.66e-05  mcm5p1f_cc_w_1_200_s_5_250 = 1.14e-12  mcm5p1f_cf_w_1_200_s_5_250 = 4.78e-11
+ mcrdlp1f_ca_w_0_150_s_0_210 = 8.27e-05  mcrdlp1f_cc_w_0_150_s_0_210 = 6.54e-11  mcrdlp1f_cf_w_0_150_s_0_210 = 8.93e-12
+ mcrdlp1f_ca_w_0_150_s_0_263 = 8.27e-05  mcrdlp1f_cc_w_0_150_s_0_263 = 5.47e-11  mcrdlp1f_cf_w_0_150_s_0_263 = 1.07e-11
+ mcrdlp1f_ca_w_0_150_s_0_315 = 8.27e-05  mcrdlp1f_cc_w_0_150_s_0_315 = 4.76e-11  mcrdlp1f_cf_w_0_150_s_0_315 = 1.24e-11
+ mcrdlp1f_ca_w_0_150_s_0_420 = 8.27e-05  mcrdlp1f_cc_w_0_150_s_0_420 = 3.73e-11  mcrdlp1f_cf_w_0_150_s_0_420 = 1.56e-11
+ mcrdlp1f_ca_w_0_150_s_0_525 = 8.27e-05  mcrdlp1f_cc_w_0_150_s_0_525 = 3.08e-11  mcrdlp1f_cf_w_0_150_s_0_525 = 1.84e-11
+ mcrdlp1f_ca_w_0_150_s_0_630 = 8.27e-05  mcrdlp1f_cc_w_0_150_s_0_630 = 2.61e-11  mcrdlp1f_cf_w_0_150_s_0_630 = 2.09e-11
+ mcrdlp1f_ca_w_0_150_s_0_840 = 8.27e-05  mcrdlp1f_cc_w_0_150_s_0_840 = 1.94e-11  mcrdlp1f_cf_w_0_150_s_0_840 = 2.52e-11
+ mcrdlp1f_ca_w_0_150_s_1_260 = 8.27e-05  mcrdlp1f_cc_w_0_150_s_1_260 = 1.14e-11  mcrdlp1f_cf_w_0_150_s_1_260 = 3.14e-11
+ mcrdlp1f_ca_w_0_150_s_2_310 = 8.27e-05  mcrdlp1f_cc_w_0_150_s_2_310 = 4.76e-12  mcrdlp1f_cf_w_0_150_s_2_310 = 3.74e-11
+ mcrdlp1f_ca_w_0_150_s_5_250 = 8.27e-05  mcrdlp1f_cc_w_0_150_s_5_250 = 9.61e-13  mcrdlp1f_cf_w_0_150_s_5_250 = 4.11e-11
+ mcrdlp1f_ca_w_1_200_s_0_210 = 8.27e-05  mcrdlp1f_cc_w_1_200_s_0_210 = 8.28e-11  mcrdlp1f_cf_w_1_200_s_0_210 = 8.87e-12
+ mcrdlp1f_ca_w_1_200_s_0_263 = 8.27e-05  mcrdlp1f_cc_w_1_200_s_0_263 = 7.09e-11  mcrdlp1f_cf_w_1_200_s_0_263 = 1.07e-11
+ mcrdlp1f_ca_w_1_200_s_0_315 = 8.27e-05  mcrdlp1f_cc_w_1_200_s_0_315 = 6.25e-11  mcrdlp1f_cf_w_1_200_s_0_315 = 1.24e-11
+ mcrdlp1f_ca_w_1_200_s_0_420 = 8.27e-05  mcrdlp1f_cc_w_1_200_s_0_420 = 5.09e-11  mcrdlp1f_cf_w_1_200_s_0_420 = 1.57e-11
+ mcrdlp1f_ca_w_1_200_s_0_525 = 8.27e-05  mcrdlp1f_cc_w_1_200_s_0_525 = 4.31e-11  mcrdlp1f_cf_w_1_200_s_0_525 = 1.86e-11
+ mcrdlp1f_ca_w_1_200_s_0_630 = 8.27e-05  mcrdlp1f_cc_w_1_200_s_0_630 = 3.74e-11  mcrdlp1f_cf_w_1_200_s_0_630 = 2.12e-11
+ mcrdlp1f_ca_w_1_200_s_0_840 = 8.27e-05  mcrdlp1f_cc_w_1_200_s_0_840 = 2.93e-11  mcrdlp1f_cf_w_1_200_s_0_840 = 2.58e-11
+ mcrdlp1f_ca_w_1_200_s_1_260 = 8.27e-05  mcrdlp1f_cc_w_1_200_s_1_260 = 1.99e-11  mcrdlp1f_cf_w_1_200_s_1_260 = 3.25e-11
+ mcrdlp1f_ca_w_1_200_s_2_310 = 8.27e-05  mcrdlp1f_cc_w_1_200_s_2_310 = 9.59e-12  mcrdlp1f_cf_w_1_200_s_2_310 = 4.13e-11
+ mcrdlp1f_ca_w_1_200_s_5_250 = 8.27e-05  mcrdlp1f_cc_w_1_200_s_5_250 = 2.47e-12  mcrdlp1f_cf_w_1_200_s_5_250 = 4.81e-11
+ mcm1l1f_ca_w_0_170_s_0_180 = 1.07e-04  mcm1l1f_cc_w_0_170_s_0_180 = 5.52e-11  mcm1l1f_cf_w_0_170_s_0_180 = 1.06e-11
+ mcm1l1f_ca_w_0_170_s_0_225 = 1.07e-04  mcm1l1f_cc_w_0_170_s_0_225 = 4.68e-11  mcm1l1f_cf_w_0_170_s_0_225 = 1.26e-11
+ mcm1l1f_ca_w_0_170_s_0_270 = 1.07e-04  mcm1l1f_cc_w_0_170_s_0_270 = 4.05e-11  mcm1l1f_cf_w_0_170_s_0_270 = 1.45e-11
+ mcm1l1f_ca_w_0_170_s_0_360 = 1.07e-04  mcm1l1f_cc_w_0_170_s_0_360 = 3.13e-11  mcm1l1f_cf_w_0_170_s_0_360 = 1.82e-11
+ mcm1l1f_ca_w_0_170_s_0_450 = 1.07e-04  mcm1l1f_cc_w_0_170_s_0_450 = 2.51e-11  mcm1l1f_cf_w_0_170_s_0_450 = 2.12e-11
+ mcm1l1f_ca_w_0_170_s_0_540 = 1.07e-04  mcm1l1f_cc_w_0_170_s_0_540 = 2.03e-11  mcm1l1f_cf_w_0_170_s_0_540 = 2.40e-11
+ mcm1l1f_ca_w_0_170_s_0_720 = 1.07e-04  mcm1l1f_cc_w_0_170_s_0_720 = 1.37e-11  mcm1l1f_cf_w_0_170_s_0_720 = 2.84e-11
+ mcm1l1f_ca_w_0_170_s_1_080 = 1.07e-04  mcm1l1f_cc_w_0_170_s_1_080 = 6.67e-12  mcm1l1f_cf_w_0_170_s_1_080 = 3.40e-11
+ mcm1l1f_ca_w_0_170_s_1_980 = 1.07e-04  mcm1l1f_cc_w_0_170_s_1_980 = 1.27e-12  mcm1l1f_cf_w_0_170_s_1_980 = 3.89e-11
+ mcm1l1f_ca_w_0_170_s_4_500 = 1.07e-04  mcm1l1f_cc_w_0_170_s_4_500 = 4.00e-14  mcm1l1f_cf_w_0_170_s_4_500 = 4.01e-11
+ mcm1l1f_ca_w_1_360_s_0_180 = 1.07e-04  mcm1l1f_cc_w_1_360_s_0_180 = 6.34e-11  mcm1l1f_cf_w_1_360_s_0_180 = 1.06e-11
+ mcm1l1f_ca_w_1_360_s_0_225 = 1.07e-04  mcm1l1f_cc_w_1_360_s_0_225 = 5.40e-11  mcm1l1f_cf_w_1_360_s_0_225 = 1.26e-11
+ mcm1l1f_ca_w_1_360_s_0_270 = 1.07e-04  mcm1l1f_cc_w_1_360_s_0_270 = 4.70e-11  mcm1l1f_cf_w_1_360_s_0_270 = 1.46e-11
+ mcm1l1f_ca_w_1_360_s_0_360 = 1.07e-04  mcm1l1f_cc_w_1_360_s_0_360 = 3.67e-11  mcm1l1f_cf_w_1_360_s_0_360 = 1.82e-11
+ mcm1l1f_ca_w_1_360_s_0_450 = 1.07e-04  mcm1l1f_cc_w_1_360_s_0_450 = 2.95e-11  mcm1l1f_cf_w_1_360_s_0_450 = 2.14e-11
+ mcm1l1f_ca_w_1_360_s_0_540 = 1.07e-04  mcm1l1f_cc_w_1_360_s_0_540 = 2.42e-11  mcm1l1f_cf_w_1_360_s_0_540 = 2.43e-11
+ mcm1l1f_ca_w_1_360_s_0_720 = 1.07e-04  mcm1l1f_cc_w_1_360_s_0_720 = 1.66e-11  mcm1l1f_cf_w_1_360_s_0_720 = 2.91e-11
+ mcm1l1f_ca_w_1_360_s_1_080 = 1.07e-04  mcm1l1f_cc_w_1_360_s_1_080 = 8.34e-12  mcm1l1f_cf_w_1_360_s_1_080 = 3.56e-11
+ mcm1l1f_ca_w_1_360_s_1_980 = 1.07e-04  mcm1l1f_cc_w_1_360_s_1_980 = 1.65e-12  mcm1l1f_cf_w_1_360_s_1_980 = 4.16e-11
+ mcm1l1f_ca_w_1_360_s_4_500 = 1.07e-04  mcm1l1f_cc_w_1_360_s_4_500 = 7.50e-14  mcm1l1f_cf_w_1_360_s_4_500 = 4.32e-11
+ mcm1l1d_ca_w_0_170_s_0_180 = 1.23e-04  mcm1l1d_cc_w_0_170_s_0_180 = 5.30e-11  mcm1l1d_cf_w_0_170_s_0_180 = 1.22e-11
+ mcm1l1d_ca_w_0_170_s_0_225 = 1.23e-04  mcm1l1d_cc_w_0_170_s_0_225 = 4.46e-11  mcm1l1d_cf_w_0_170_s_0_225 = 1.45e-11
+ mcm1l1d_ca_w_0_170_s_0_270 = 1.23e-04  mcm1l1d_cc_w_0_170_s_0_270 = 3.81e-11  mcm1l1d_cf_w_0_170_s_0_270 = 1.66e-11
+ mcm1l1d_ca_w_0_170_s_0_360 = 1.23e-04  mcm1l1d_cc_w_0_170_s_0_360 = 2.88e-11  mcm1l1d_cf_w_0_170_s_0_360 = 2.06e-11
+ mcm1l1d_ca_w_0_170_s_0_450 = 1.23e-04  mcm1l1d_cc_w_0_170_s_0_450 = 2.24e-11  mcm1l1d_cf_w_0_170_s_0_450 = 2.39e-11
+ mcm1l1d_ca_w_0_170_s_0_540 = 1.23e-04  mcm1l1d_cc_w_0_170_s_0_540 = 1.77e-11  mcm1l1d_cf_w_0_170_s_0_540 = 2.69e-11
+ mcm1l1d_ca_w_0_170_s_0_720 = 1.23e-04  mcm1l1d_cc_w_0_170_s_0_720 = 1.13e-11  mcm1l1d_cf_w_0_170_s_0_720 = 3.14e-11
+ mcm1l1d_ca_w_0_170_s_1_080 = 1.23e-04  mcm1l1d_cc_w_0_170_s_1_080 = 4.82e-12  mcm1l1d_cf_w_0_170_s_1_080 = 3.68e-11
+ mcm1l1d_ca_w_0_170_s_1_980 = 1.23e-04  mcm1l1d_cc_w_0_170_s_1_980 = 6.45e-13  mcm1l1d_cf_w_0_170_s_1_980 = 4.07e-11
+ mcm1l1d_ca_w_0_170_s_4_500 = 1.23e-04  mcm1l1d_cc_w_0_170_s_4_500 = 2.00e-14  mcm1l1d_cf_w_0_170_s_4_500 = 4.13e-11
+ mcm1l1d_ca_w_1_360_s_0_180 = 1.23e-04  mcm1l1d_cc_w_1_360_s_0_180 = 5.91e-11  mcm1l1d_cf_w_1_360_s_0_180 = 1.21e-11
+ mcm1l1d_ca_w_1_360_s_0_225 = 1.23e-04  mcm1l1d_cc_w_1_360_s_0_225 = 4.98e-11  mcm1l1d_cf_w_1_360_s_0_225 = 1.44e-11
+ mcm1l1d_ca_w_1_360_s_0_270 = 1.23e-04  mcm1l1d_cc_w_1_360_s_0_270 = 4.26e-11  mcm1l1d_cf_w_1_360_s_0_270 = 1.66e-11
+ mcm1l1d_ca_w_1_360_s_0_360 = 1.23e-04  mcm1l1d_cc_w_1_360_s_0_360 = 3.25e-11  mcm1l1d_cf_w_1_360_s_0_360 = 2.06e-11
+ mcm1l1d_ca_w_1_360_s_0_450 = 1.23e-04  mcm1l1d_cc_w_1_360_s_0_450 = 2.53e-11  mcm1l1d_cf_w_1_360_s_0_450 = 2.42e-11
+ mcm1l1d_ca_w_1_360_s_0_540 = 1.23e-04  mcm1l1d_cc_w_1_360_s_0_540 = 2.00e-11  mcm1l1d_cf_w_1_360_s_0_540 = 2.73e-11
+ mcm1l1d_ca_w_1_360_s_0_720 = 1.23e-04  mcm1l1d_cc_w_1_360_s_0_720 = 1.30e-11  mcm1l1d_cf_w_1_360_s_0_720 = 3.22e-11
+ mcm1l1d_ca_w_1_360_s_1_080 = 1.23e-04  mcm1l1d_cc_w_1_360_s_1_080 = 5.60e-12  mcm1l1d_cf_w_1_360_s_1_080 = 3.82e-11
+ mcm1l1d_ca_w_1_360_s_1_980 = 1.23e-04  mcm1l1d_cc_w_1_360_s_1_980 = 7.85e-13  mcm1l1d_cf_w_1_360_s_1_980 = 4.27e-11
+ mcm1l1d_ca_w_1_360_s_4_500 = 1.23e-04  mcm1l1d_cc_w_1_360_s_4_500 = 5.00e-14  mcm1l1d_cf_w_1_360_s_4_500 = 4.35e-11
+ mcm1l1p1_ca_w_0_170_s_0_180 = 1.42e-04  mcm1l1p1_cc_w_0_170_s_0_180 = 5.07e-11  mcm1l1p1_cf_w_0_170_s_0_180 = 1.40e-11
+ mcm1l1p1_ca_w_0_170_s_0_225 = 1.42e-04  mcm1l1p1_cc_w_0_170_s_0_225 = 4.21e-11  mcm1l1p1_cf_w_0_170_s_0_225 = 1.66e-11
+ mcm1l1p1_ca_w_0_170_s_0_270 = 1.42e-04  mcm1l1p1_cc_w_0_170_s_0_270 = 3.56e-11  mcm1l1p1_cf_w_0_170_s_0_270 = 1.90e-11
+ mcm1l1p1_ca_w_0_170_s_0_360 = 1.42e-04  mcm1l1p1_cc_w_0_170_s_0_360 = 2.62e-11  mcm1l1p1_cf_w_0_170_s_0_360 = 2.34e-11
+ mcm1l1p1_ca_w_0_170_s_0_450 = 1.42e-04  mcm1l1p1_cc_w_0_170_s_0_450 = 1.99e-11  mcm1l1p1_cf_w_0_170_s_0_450 = 2.70e-11
+ mcm1l1p1_ca_w_0_170_s_0_540 = 1.42e-04  mcm1l1p1_cc_w_0_170_s_0_540 = 1.52e-11  mcm1l1p1_cf_w_0_170_s_0_540 = 3.01e-11
+ mcm1l1p1_ca_w_0_170_s_0_720 = 1.42e-04  mcm1l1p1_cc_w_0_170_s_0_720 = 9.16e-12  mcm1l1p1_cf_w_0_170_s_0_720 = 3.47e-11
+ mcm1l1p1_ca_w_0_170_s_1_080 = 1.42e-04  mcm1l1p1_cc_w_0_170_s_1_080 = 3.42e-12  mcm1l1p1_cf_w_0_170_s_1_080 = 3.97e-11
+ mcm1l1p1_ca_w_0_170_s_1_980 = 1.42e-04  mcm1l1p1_cc_w_0_170_s_1_980 = 3.45e-13  mcm1l1p1_cf_w_0_170_s_1_980 = 4.26e-11
+ mcm1l1p1_ca_w_0_170_s_4_500 = 1.42e-04  mcm1l1p1_cc_w_0_170_s_4_500 = 2.50e-14  mcm1l1p1_cf_w_0_170_s_4_500 = 4.29e-11
+ mcm1l1p1_ca_w_1_360_s_0_180 = 1.42e-04  mcm1l1p1_cc_w_1_360_s_0_180 = 5.49e-11  mcm1l1p1_cf_w_1_360_s_0_180 = 1.39e-11
+ mcm1l1p1_ca_w_1_360_s_0_225 = 1.42e-04  mcm1l1p1_cc_w_1_360_s_0_225 = 4.57e-11  mcm1l1p1_cf_w_1_360_s_0_225 = 1.65e-11
+ mcm1l1p1_ca_w_1_360_s_0_270 = 1.42e-04  mcm1l1p1_cc_w_1_360_s_0_270 = 3.87e-11  mcm1l1p1_cf_w_1_360_s_0_270 = 1.90e-11
+ mcm1l1p1_ca_w_1_360_s_0_360 = 1.42e-04  mcm1l1p1_cc_w_1_360_s_0_360 = 2.85e-11  mcm1l1p1_cf_w_1_360_s_0_360 = 2.35e-11
+ mcm1l1p1_ca_w_1_360_s_0_450 = 1.42e-04  mcm1l1p1_cc_w_1_360_s_0_450 = 2.17e-11  mcm1l1p1_cf_w_1_360_s_0_450 = 2.73e-11
+ mcm1l1p1_ca_w_1_360_s_0_540 = 1.42e-04  mcm1l1p1_cc_w_1_360_s_0_540 = 1.67e-11  mcm1l1p1_cf_w_1_360_s_0_540 = 3.05e-11
+ mcm1l1p1_ca_w_1_360_s_0_720 = 1.42e-04  mcm1l1p1_cc_w_1_360_s_0_720 = 1.01e-11  mcm1l1p1_cf_w_1_360_s_0_720 = 3.54e-11
+ mcm1l1p1_ca_w_1_360_s_1_080 = 1.42e-04  mcm1l1p1_cc_w_1_360_s_1_080 = 3.85e-12  mcm1l1p1_cf_w_1_360_s_1_080 = 4.08e-11
+ mcm1l1p1_ca_w_1_360_s_1_980 = 1.42e-04  mcm1l1p1_cc_w_1_360_s_1_980 = 3.50e-13  mcm1l1p1_cf_w_1_360_s_1_980 = 4.41e-11
+ mcm1l1p1_ca_w_1_360_s_4_500 = 1.42e-04  mcm1l1p1_cc_w_1_360_s_4_500 = 5.00e-14  mcm1l1p1_cf_w_1_360_s_4_500 = 4.44e-11
+ mcm2l1f_ca_w_0_170_s_0_180 = 5.80e-05  mcm2l1f_cc_w_0_170_s_0_180 = 6.11e-11  mcm2l1f_cf_w_0_170_s_0_180 = 6.02e-12
+ mcm2l1f_ca_w_0_170_s_0_225 = 5.80e-05  mcm2l1f_cc_w_0_170_s_0_225 = 5.30e-11  mcm2l1f_cf_w_0_170_s_0_225 = 7.21e-12
+ mcm2l1f_ca_w_0_170_s_0_270 = 5.80e-05  mcm2l1f_cc_w_0_170_s_0_270 = 4.72e-11  mcm2l1f_cf_w_0_170_s_0_270 = 8.35e-12
+ mcm2l1f_ca_w_0_170_s_0_360 = 5.80e-05  mcm2l1f_cc_w_0_170_s_0_360 = 3.84e-11  mcm2l1f_cf_w_0_170_s_0_360 = 1.07e-11
+ mcm2l1f_ca_w_0_170_s_0_450 = 5.80e-05  mcm2l1f_cc_w_0_170_s_0_450 = 3.24e-11  mcm2l1f_cf_w_0_170_s_0_450 = 1.27e-11
+ mcm2l1f_ca_w_0_170_s_0_540 = 5.80e-05  mcm2l1f_cc_w_0_170_s_0_540 = 2.75e-11  mcm2l1f_cf_w_0_170_s_0_540 = 1.47e-11
+ mcm2l1f_ca_w_0_170_s_0_720 = 5.80e-05  mcm2l1f_cc_w_0_170_s_0_720 = 2.08e-11  mcm2l1f_cf_w_0_170_s_0_720 = 1.81e-11
+ mcm2l1f_ca_w_0_170_s_1_080 = 5.80e-05  mcm2l1f_cc_w_0_170_s_1_080 = 1.25e-11  mcm2l1f_cf_w_0_170_s_1_080 = 2.34e-11
+ mcm2l1f_ca_w_0_170_s_1_980 = 5.80e-05  mcm2l1f_cc_w_0_170_s_1_980 = 3.94e-12  mcm2l1f_cf_w_0_170_s_1_980 = 3.03e-11
+ mcm2l1f_ca_w_0_170_s_4_500 = 5.80e-05  mcm2l1f_cc_w_0_170_s_4_500 = 2.10e-13  mcm2l1f_cf_w_0_170_s_4_500 = 3.38e-11
+ mcm2l1f_ca_w_1_360_s_0_180 = 5.80e-05  mcm2l1f_cc_w_1_360_s_0_180 = 7.39e-11  mcm2l1f_cf_w_1_360_s_0_180 = 5.99e-12
+ mcm2l1f_ca_w_1_360_s_0_225 = 5.80e-05  mcm2l1f_cc_w_1_360_s_0_225 = 6.46e-11  mcm2l1f_cf_w_1_360_s_0_225 = 7.20e-12
+ mcm2l1f_ca_w_1_360_s_0_270 = 5.80e-05  mcm2l1f_cc_w_1_360_s_0_270 = 5.75e-11  mcm2l1f_cf_w_1_360_s_0_270 = 8.38e-12
+ mcm2l1f_ca_w_1_360_s_0_360 = 5.80e-05  mcm2l1f_cc_w_1_360_s_0_360 = 4.71e-11  mcm2l1f_cf_w_1_360_s_0_360 = 1.07e-11
+ mcm2l1f_ca_w_1_360_s_0_450 = 5.80e-05  mcm2l1f_cc_w_1_360_s_0_450 = 3.97e-11  mcm2l1f_cf_w_1_360_s_0_450 = 1.28e-11
+ mcm2l1f_ca_w_1_360_s_0_540 = 5.80e-05  mcm2l1f_cc_w_1_360_s_0_540 = 3.40e-11  mcm2l1f_cf_w_1_360_s_0_540 = 1.49e-11
+ mcm2l1f_ca_w_1_360_s_0_720 = 5.80e-05  mcm2l1f_cc_w_1_360_s_0_720 = 2.58e-11  mcm2l1f_cf_w_1_360_s_0_720 = 1.85e-11
+ mcm2l1f_ca_w_1_360_s_1_080 = 5.80e-05  mcm2l1f_cc_w_1_360_s_1_080 = 1.57e-11  mcm2l1f_cf_w_1_360_s_1_080 = 2.44e-11
+ mcm2l1f_ca_w_1_360_s_1_980 = 5.80e-05  mcm2l1f_cc_w_1_360_s_1_980 = 5.08e-12  mcm2l1f_cf_w_1_360_s_1_980 = 3.28e-11
+ mcm2l1f_ca_w_1_360_s_4_500 = 5.80e-05  mcm2l1f_cc_w_1_360_s_4_500 = 2.80e-13  mcm2l1f_cf_w_1_360_s_4_500 = 3.73e-11
+ mcm2l1d_ca_w_0_170_s_0_180 = 7.39e-05  mcm2l1d_cc_w_0_170_s_0_180 = 5.90e-11  mcm2l1d_cf_w_0_170_s_0_180 = 7.61e-12
+ mcm2l1d_ca_w_0_170_s_0_225 = 7.39e-05  mcm2l1d_cc_w_0_170_s_0_225 = 5.08e-11  mcm2l1d_cf_w_0_170_s_0_225 = 9.10e-12
+ mcm2l1d_ca_w_0_170_s_0_270 = 7.39e-05  mcm2l1d_cc_w_0_170_s_0_270 = 4.47e-11  mcm2l1d_cf_w_0_170_s_0_270 = 1.05e-11
+ mcm2l1d_ca_w_0_170_s_0_360 = 7.39e-05  mcm2l1d_cc_w_0_170_s_0_360 = 3.56e-11  mcm2l1d_cf_w_0_170_s_0_360 = 1.34e-11
+ mcm2l1d_ca_w_0_170_s_0_450 = 7.39e-05  mcm2l1d_cc_w_0_170_s_0_450 = 2.95e-11  mcm2l1d_cf_w_0_170_s_0_450 = 1.58e-11
+ mcm2l1d_ca_w_0_170_s_0_540 = 7.39e-05  mcm2l1d_cc_w_0_170_s_0_540 = 2.46e-11  mcm2l1d_cf_w_0_170_s_0_540 = 1.81e-11
+ mcm2l1d_ca_w_0_170_s_0_720 = 7.39e-05  mcm2l1d_cc_w_0_170_s_0_720 = 1.78e-11  mcm2l1d_cf_w_0_170_s_0_720 = 2.20e-11
+ mcm2l1d_ca_w_0_170_s_1_080 = 7.39e-05  mcm2l1d_cc_w_0_170_s_1_080 = 9.83e-12  mcm2l1d_cf_w_0_170_s_1_080 = 2.76e-11
+ mcm2l1d_ca_w_0_170_s_1_980 = 7.39e-05  mcm2l1d_cc_w_0_170_s_1_980 = 2.47e-12  mcm2l1d_cf_w_0_170_s_1_980 = 3.39e-11
+ mcm2l1d_ca_w_0_170_s_4_500 = 7.39e-05  mcm2l1d_cc_w_0_170_s_4_500 = 9.50e-14  mcm2l1d_cf_w_0_170_s_4_500 = 3.62e-11
+ mcm2l1d_ca_w_1_360_s_0_180 = 7.39e-05  mcm2l1d_cc_w_1_360_s_0_180 = 6.93e-11  mcm2l1d_cf_w_1_360_s_0_180 = 7.59e-12
+ mcm2l1d_ca_w_1_360_s_0_225 = 7.39e-05  mcm2l1d_cc_w_1_360_s_0_225 = 6.00e-11  mcm2l1d_cf_w_1_360_s_0_225 = 9.09e-12
+ mcm2l1d_ca_w_1_360_s_0_270 = 7.39e-05  mcm2l1d_cc_w_1_360_s_0_270 = 5.28e-11  mcm2l1d_cf_w_1_360_s_0_270 = 1.06e-11
+ mcm2l1d_ca_w_1_360_s_0_360 = 7.39e-05  mcm2l1d_cc_w_1_360_s_0_360 = 4.25e-11  mcm2l1d_cf_w_1_360_s_0_360 = 1.33e-11
+ mcm2l1d_ca_w_1_360_s_0_450 = 7.39e-05  mcm2l1d_cc_w_1_360_s_0_450 = 3.52e-11  mcm2l1d_cf_w_1_360_s_0_450 = 1.60e-11
+ mcm2l1d_ca_w_1_360_s_0_540 = 7.39e-05  mcm2l1d_cc_w_1_360_s_0_540 = 2.96e-11  mcm2l1d_cf_w_1_360_s_0_540 = 1.83e-11
+ mcm2l1d_ca_w_1_360_s_0_720 = 7.39e-05  mcm2l1d_cc_w_1_360_s_0_720 = 2.16e-11  mcm2l1d_cf_w_1_360_s_0_720 = 2.26e-11
+ mcm2l1d_ca_w_1_360_s_1_080 = 7.39e-05  mcm2l1d_cc_w_1_360_s_1_080 = 1.21e-11  mcm2l1d_cf_w_1_360_s_1_080 = 2.89e-11
+ mcm2l1d_ca_w_1_360_s_1_980 = 7.39e-05  mcm2l1d_cc_w_1_360_s_1_980 = 3.16e-12  mcm2l1d_cf_w_1_360_s_1_980 = 3.65e-11
+ mcm2l1d_ca_w_1_360_s_4_500 = 7.39e-05  mcm2l1d_cc_w_1_360_s_4_500 = 1.50e-13  mcm2l1d_cf_w_1_360_s_4_500 = 3.94e-11
+ mcm2l1p1_ca_w_0_170_s_0_180 = 9.32e-05  mcm2l1p1_cc_w_0_170_s_0_180 = 5.66e-11  mcm2l1p1_cf_w_0_170_s_0_180 = 9.50e-12
+ mcm2l1p1_ca_w_0_170_s_0_225 = 9.32e-05  mcm2l1p1_cc_w_0_170_s_0_225 = 4.83e-11  mcm2l1p1_cf_w_0_170_s_0_225 = 1.13e-11
+ mcm2l1p1_ca_w_0_170_s_0_270 = 9.32e-05  mcm2l1p1_cc_w_0_170_s_0_270 = 4.20e-11  mcm2l1p1_cf_w_0_170_s_0_270 = 1.30e-11
+ mcm2l1p1_ca_w_0_170_s_0_360 = 9.32e-05  mcm2l1p1_cc_w_0_170_s_0_360 = 3.29e-11  mcm2l1p1_cf_w_0_170_s_0_360 = 1.64e-11
+ mcm2l1p1_ca_w_0_170_s_0_450 = 9.32e-05  mcm2l1p1_cc_w_0_170_s_0_450 = 2.66e-11  mcm2l1p1_cf_w_0_170_s_0_450 = 1.92e-11
+ mcm2l1p1_ca_w_0_170_s_0_540 = 9.32e-05  mcm2l1p1_cc_w_0_170_s_0_540 = 2.18e-11  mcm2l1p1_cf_w_0_170_s_0_540 = 2.19e-11
+ mcm2l1p1_ca_w_0_170_s_0_720 = 9.32e-05  mcm2l1p1_cc_w_0_170_s_0_720 = 1.51e-11  mcm2l1p1_cf_w_0_170_s_0_720 = 2.62e-11
+ mcm2l1p1_ca_w_0_170_s_1_080 = 9.32e-05  mcm2l1p1_cc_w_0_170_s_1_080 = 7.66e-12  mcm2l1p1_cf_w_0_170_s_1_080 = 3.19e-11
+ mcm2l1p1_ca_w_0_170_s_1_980 = 9.32e-05  mcm2l1p1_cc_w_0_170_s_1_980 = 1.61e-12  mcm2l1p1_cf_w_0_170_s_1_980 = 3.73e-11
+ mcm2l1p1_ca_w_0_170_s_4_500 = 9.32e-05  mcm2l1p1_cc_w_0_170_s_4_500 = 5.00e-14  mcm2l1p1_cf_w_0_170_s_4_500 = 3.88e-11
+ mcm2l1p1_ca_w_1_360_s_0_180 = 9.32e-05  mcm2l1p1_cc_w_1_360_s_0_180 = 6.53e-11  mcm2l1p1_cf_w_1_360_s_0_180 = 9.47e-12
+ mcm2l1p1_ca_w_1_360_s_0_225 = 9.32e-05  mcm2l1p1_cc_w_1_360_s_0_225 = 5.60e-11  mcm2l1p1_cf_w_1_360_s_0_225 = 1.13e-11
+ mcm2l1p1_ca_w_1_360_s_0_270 = 9.32e-05  mcm2l1p1_cc_w_1_360_s_0_270 = 4.90e-11  mcm2l1p1_cf_w_1_360_s_0_270 = 1.31e-11
+ mcm2l1p1_ca_w_1_360_s_0_360 = 9.32e-05  mcm2l1p1_cc_w_1_360_s_0_360 = 3.87e-11  mcm2l1p1_cf_w_1_360_s_0_360 = 1.64e-11
+ mcm2l1p1_ca_w_1_360_s_0_450 = 9.32e-05  mcm2l1p1_cc_w_1_360_s_0_450 = 3.14e-11  mcm2l1p1_cf_w_1_360_s_0_450 = 1.95e-11
+ mcm2l1p1_ca_w_1_360_s_0_540 = 9.32e-05  mcm2l1p1_cc_w_1_360_s_0_540 = 2.60e-11  mcm2l1p1_cf_w_1_360_s_0_540 = 2.22e-11
+ mcm2l1p1_ca_w_1_360_s_0_720 = 9.32e-05  mcm2l1p1_cc_w_1_360_s_0_720 = 1.82e-11  mcm2l1p1_cf_w_1_360_s_0_720 = 2.69e-11
+ mcm2l1p1_ca_w_1_360_s_1_080 = 9.32e-05  mcm2l1p1_cc_w_1_360_s_1_080 = 9.53e-12  mcm2l1p1_cf_w_1_360_s_1_080 = 3.33e-11
+ mcm2l1p1_ca_w_1_360_s_1_980 = 9.32e-05  mcm2l1p1_cc_w_1_360_s_1_980 = 2.06e-12  mcm2l1p1_cf_w_1_360_s_1_980 = 4.00e-11
+ mcm2l1p1_ca_w_1_360_s_4_500 = 9.32e-05  mcm2l1p1_cc_w_1_360_s_4_500 = 2.50e-14  mcm2l1p1_cf_w_1_360_s_4_500 = 4.20e-11
+ mcm3l1f_ca_w_0_170_s_0_180 = 4.57e-05  mcm3l1f_cc_w_0_170_s_0_180 = 6.29e-11  mcm3l1f_cf_w_0_170_s_0_180 = 4.78e-12
+ mcm3l1f_ca_w_0_170_s_0_225 = 4.57e-05  mcm3l1f_cc_w_0_170_s_0_225 = 5.49e-11  mcm3l1f_cf_w_0_170_s_0_225 = 5.73e-12
+ mcm3l1f_ca_w_0_170_s_0_270 = 4.57e-05  mcm3l1f_cc_w_0_170_s_0_270 = 4.94e-11  mcm3l1f_cf_w_0_170_s_0_270 = 6.65e-12
+ mcm3l1f_ca_w_0_170_s_0_360 = 4.57e-05  mcm3l1f_cc_w_0_170_s_0_360 = 4.07e-11  mcm3l1f_cf_w_0_170_s_0_360 = 8.65e-12
+ mcm3l1f_ca_w_0_170_s_0_450 = 4.57e-05  mcm3l1f_cc_w_0_170_s_0_450 = 3.50e-11  mcm3l1f_cf_w_0_170_s_0_450 = 1.02e-11
+ mcm3l1f_ca_w_0_170_s_0_540 = 4.57e-05  mcm3l1f_cc_w_0_170_s_0_540 = 3.03e-11  mcm3l1f_cf_w_0_170_s_0_540 = 1.20e-11
+ mcm3l1f_ca_w_0_170_s_0_720 = 4.57e-05  mcm3l1f_cc_w_0_170_s_0_720 = 2.37e-11  mcm3l1f_cf_w_0_170_s_0_720 = 1.49e-11
+ mcm3l1f_ca_w_0_170_s_1_080 = 4.57e-05  mcm3l1f_cc_w_0_170_s_1_080 = 1.55e-11  mcm3l1f_cf_w_0_170_s_1_080 = 1.96e-11
+ mcm3l1f_ca_w_0_170_s_1_980 = 4.57e-05  mcm3l1f_cc_w_0_170_s_1_980 = 6.09e-12  mcm3l1f_cf_w_0_170_s_1_980 = 2.67e-11
+ mcm3l1f_ca_w_0_170_s_4_500 = 4.57e-05  mcm3l1f_cc_w_0_170_s_4_500 = 5.95e-13  mcm3l1f_cf_w_0_170_s_4_500 = 3.17e-11
+ mcm3l1f_ca_w_1_360_s_0_180 = 4.57e-05  mcm3l1f_cc_w_1_360_s_0_180 = 7.91e-11  mcm3l1f_cf_w_1_360_s_0_180 = 4.75e-12
+ mcm3l1f_ca_w_1_360_s_0_225 = 4.57e-05  mcm3l1f_cc_w_1_360_s_0_225 = 6.98e-11  mcm3l1f_cf_w_1_360_s_0_225 = 5.72e-12
+ mcm3l1f_ca_w_1_360_s_0_270 = 4.57e-05  mcm3l1f_cc_w_1_360_s_0_270 = 6.27e-11  mcm3l1f_cf_w_1_360_s_0_270 = 6.67e-12
+ mcm3l1f_ca_w_1_360_s_0_360 = 4.57e-05  mcm3l1f_cc_w_1_360_s_0_360 = 5.24e-11  mcm3l1f_cf_w_1_360_s_0_360 = 8.52e-12
+ mcm3l1f_ca_w_1_360_s_0_450 = 4.57e-05  mcm3l1f_cc_w_1_360_s_0_450 = 4.50e-11  mcm3l1f_cf_w_1_360_s_0_450 = 1.03e-11
+ mcm3l1f_ca_w_1_360_s_0_540 = 4.57e-05  mcm3l1f_cc_w_1_360_s_0_540 = 3.93e-11  mcm3l1f_cf_w_1_360_s_0_540 = 1.20e-11
+ mcm3l1f_ca_w_1_360_s_0_720 = 4.57e-05  mcm3l1f_cc_w_1_360_s_0_720 = 3.10e-11  mcm3l1f_cf_w_1_360_s_0_720 = 1.51e-11
+ mcm3l1f_ca_w_1_360_s_1_080 = 4.57e-05  mcm3l1f_cc_w_1_360_s_1_080 = 2.06e-11  mcm3l1f_cf_w_1_360_s_1_080 = 2.05e-11
+ mcm3l1f_ca_w_1_360_s_1_980 = 4.57e-05  mcm3l1f_cc_w_1_360_s_1_980 = 8.43e-12  mcm3l1f_cf_w_1_360_s_1_980 = 2.91e-11
+ mcm3l1f_ca_w_1_360_s_4_500 = 4.57e-05  mcm3l1f_cc_w_1_360_s_4_500 = 8.60e-13  mcm3l1f_cf_w_1_360_s_4_500 = 3.60e-11
+ mcm3l1d_ca_w_0_170_s_0_180 = 6.16e-05  mcm3l1d_cc_w_0_170_s_0_180 = 6.07e-11  mcm3l1d_cf_w_0_170_s_0_180 = 6.38e-12
+ mcm3l1d_ca_w_0_170_s_0_225 = 6.16e-05  mcm3l1d_cc_w_0_170_s_0_225 = 5.26e-11  mcm3l1d_cf_w_0_170_s_0_225 = 7.64e-12
+ mcm3l1d_ca_w_0_170_s_0_270 = 6.16e-05  mcm3l1d_cc_w_0_170_s_0_270 = 4.69e-11  mcm3l1d_cf_w_0_170_s_0_270 = 8.84e-12
+ mcm3l1d_ca_w_0_170_s_0_360 = 6.16e-05  mcm3l1d_cc_w_0_170_s_0_360 = 3.79e-11  mcm3l1d_cf_w_0_170_s_0_360 = 1.14e-11
+ mcm3l1d_ca_w_0_170_s_0_450 = 6.16e-05  mcm3l1d_cc_w_0_170_s_0_450 = 3.21e-11  mcm3l1d_cf_w_0_170_s_0_450 = 1.34e-11
+ mcm3l1d_ca_w_0_170_s_0_540 = 6.16e-05  mcm3l1d_cc_w_0_170_s_0_540 = 2.72e-11  mcm3l1d_cf_w_0_170_s_0_540 = 1.55e-11
+ mcm3l1d_ca_w_0_170_s_0_720 = 6.16e-05  mcm3l1d_cc_w_0_170_s_0_720 = 2.05e-11  mcm3l1d_cf_w_0_170_s_0_720 = 1.91e-11
+ mcm3l1d_ca_w_0_170_s_1_080 = 6.16e-05  mcm3l1d_cc_w_0_170_s_1_080 = 1.24e-11  mcm3l1d_cf_w_0_170_s_1_080 = 2.44e-11
+ mcm3l1d_ca_w_0_170_s_1_980 = 6.16e-05  mcm3l1d_cc_w_0_170_s_1_980 = 4.14e-12  mcm3l1d_cf_w_0_170_s_1_980 = 3.12e-11
+ mcm3l1d_ca_w_0_170_s_4_500 = 6.16e-05  mcm3l1d_cc_w_0_170_s_4_500 = 2.95e-13  mcm3l1d_cf_w_0_170_s_4_500 = 3.48e-11
+ mcm3l1d_ca_w_1_360_s_0_180 = 6.16e-05  mcm3l1d_cc_w_1_360_s_0_180 = 7.44e-11  mcm3l1d_cf_w_1_360_s_0_180 = 6.36e-12
+ mcm3l1d_ca_w_1_360_s_0_225 = 6.16e-05  mcm3l1d_cc_w_1_360_s_0_225 = 6.52e-11  mcm3l1d_cf_w_1_360_s_0_225 = 7.63e-12
+ mcm3l1d_ca_w_1_360_s_0_270 = 6.16e-05  mcm3l1d_cc_w_1_360_s_0_270 = 5.81e-11  mcm3l1d_cf_w_1_360_s_0_270 = 8.88e-12
+ mcm3l1d_ca_w_1_360_s_0_360 = 6.16e-05  mcm3l1d_cc_w_1_360_s_0_360 = 4.77e-11  mcm3l1d_cf_w_1_360_s_0_360 = 1.13e-11
+ mcm3l1d_ca_w_1_360_s_0_450 = 6.16e-05  mcm3l1d_cc_w_1_360_s_0_450 = 4.04e-11  mcm3l1d_cf_w_1_360_s_0_450 = 1.35e-11
+ mcm3l1d_ca_w_1_360_s_0_540 = 6.16e-05  mcm3l1d_cc_w_1_360_s_0_540 = 3.48e-11  mcm3l1d_cf_w_1_360_s_0_540 = 1.56e-11
+ mcm3l1d_ca_w_1_360_s_0_720 = 6.16e-05  mcm3l1d_cc_w_1_360_s_0_720 = 2.66e-11  mcm3l1d_cf_w_1_360_s_0_720 = 1.94e-11
+ mcm3l1d_ca_w_1_360_s_1_080 = 6.16e-05  mcm3l1d_cc_w_1_360_s_1_080 = 1.67e-11  mcm3l1d_cf_w_1_360_s_1_080 = 2.55e-11
+ mcm3l1d_ca_w_1_360_s_1_980 = 6.16e-05  mcm3l1d_cc_w_1_360_s_1_980 = 5.91e-12  mcm3l1d_cf_w_1_360_s_1_980 = 3.40e-11
+ mcm3l1d_ca_w_1_360_s_4_500 = 6.16e-05  mcm3l1d_cc_w_1_360_s_4_500 = 4.40e-13  mcm3l1d_cf_w_1_360_s_4_500 = 3.92e-11
+ mcm3l1p1_ca_w_0_170_s_0_180 = 8.09e-05  mcm3l1p1_cc_w_0_170_s_0_180 = 5.83e-11  mcm3l1p1_cf_w_0_170_s_0_180 = 8.28e-12
+ mcm3l1p1_ca_w_0_170_s_0_225 = 8.09e-05  mcm3l1p1_cc_w_0_170_s_0_225 = 5.00e-11  mcm3l1p1_cf_w_0_170_s_0_225 = 9.88e-12
+ mcm3l1p1_ca_w_0_170_s_0_270 = 8.09e-05  mcm3l1p1_cc_w_0_170_s_0_270 = 4.42e-11  mcm3l1p1_cf_w_0_170_s_0_270 = 1.14e-11
+ mcm3l1p1_ca_w_0_170_s_0_360 = 8.09e-05  mcm3l1p1_cc_w_0_170_s_0_360 = 3.51e-11  mcm3l1p1_cf_w_0_170_s_0_360 = 1.45e-11
+ mcm3l1p1_ca_w_0_170_s_0_450 = 8.09e-05  mcm3l1p1_cc_w_0_170_s_0_450 = 2.91e-11  mcm3l1p1_cf_w_0_170_s_0_450 = 1.70e-11
+ mcm3l1p1_ca_w_0_170_s_0_540 = 8.09e-05  mcm3l1p1_cc_w_0_170_s_0_540 = 2.42e-11  mcm3l1p1_cf_w_0_170_s_0_540 = 1.95e-11
+ mcm3l1p1_ca_w_0_170_s_0_720 = 8.09e-05  mcm3l1p1_cc_w_0_170_s_0_720 = 1.76e-11  mcm3l1p1_cf_w_0_170_s_0_720 = 2.35e-11
+ mcm3l1p1_ca_w_0_170_s_1_080 = 8.09e-05  mcm3l1p1_cc_w_0_170_s_1_080 = 9.91e-12  mcm3l1p1_cf_w_0_170_s_1_080 = 2.91e-11
+ mcm3l1p1_ca_w_0_170_s_1_980 = 8.09e-05  mcm3l1p1_cc_w_0_170_s_1_980 = 2.87e-12  mcm3l1p1_cf_w_0_170_s_1_980 = 3.53e-11
+ mcm3l1p1_ca_w_0_170_s_4_500 = 8.09e-05  mcm3l1p1_cc_w_0_170_s_4_500 = 1.80e-13  mcm3l1p1_cf_w_0_170_s_4_500 = 3.79e-11
+ mcm3l1p1_ca_w_1_360_s_0_180 = 8.09e-05  mcm3l1p1_cc_w_1_360_s_0_180 = 7.05e-11  mcm3l1p1_cf_w_1_360_s_0_180 = 8.29e-12
+ mcm3l1p1_ca_w_1_360_s_0_225 = 8.09e-05  mcm3l1p1_cc_w_1_360_s_0_225 = 6.13e-11  mcm3l1p1_cf_w_1_360_s_0_225 = 9.92e-12
+ mcm3l1p1_ca_w_1_360_s_0_270 = 8.09e-05  mcm3l1p1_cc_w_1_360_s_0_270 = 5.42e-11  mcm3l1p1_cf_w_1_360_s_0_270 = 1.15e-11
+ mcm3l1p1_ca_w_1_360_s_0_360 = 8.09e-05  mcm3l1p1_cc_w_1_360_s_0_360 = 4.40e-11  mcm3l1p1_cf_w_1_360_s_0_360 = 1.44e-11
+ mcm3l1p1_ca_w_1_360_s_0_450 = 8.09e-05  mcm3l1p1_cc_w_1_360_s_0_450 = 3.66e-11  mcm3l1p1_cf_w_1_360_s_0_450 = 1.72e-11
+ mcm3l1p1_ca_w_1_360_s_0_540 = 8.09e-05  mcm3l1p1_cc_w_1_360_s_0_540 = 3.11e-11  mcm3l1p1_cf_w_1_360_s_0_540 = 1.97e-11
+ mcm3l1p1_ca_w_1_360_s_0_720 = 8.09e-05  mcm3l1p1_cc_w_1_360_s_0_720 = 2.32e-11  mcm3l1p1_cf_w_1_360_s_0_720 = 2.41e-11
+ mcm3l1p1_ca_w_1_360_s_1_080 = 8.09e-05  mcm3l1p1_cc_w_1_360_s_1_080 = 1.38e-11  mcm3l1p1_cf_w_1_360_s_1_080 = 3.06e-11
+ mcm3l1p1_ca_w_1_360_s_1_980 = 8.09e-05  mcm3l1p1_cc_w_1_360_s_1_980 = 4.41e-12  mcm3l1p1_cf_w_1_360_s_1_980 = 3.86e-11
+ mcm3l1p1_ca_w_1_360_s_4_500 = 8.09e-05  mcm3l1p1_cc_w_1_360_s_4_500 = 2.50e-13  mcm3l1p1_cf_w_1_360_s_4_500 = 4.25e-11
+ mcm4l1f_ca_w_0_170_s_0_180 = 3.93e-05  mcm4l1f_cc_w_0_170_s_0_180 = 6.38e-11  mcm4l1f_cf_w_0_170_s_0_180 = 4.12e-12
+ mcm4l1f_ca_w_0_170_s_0_225 = 3.93e-05  mcm4l1f_cc_w_0_170_s_0_225 = 5.59e-11  mcm4l1f_cf_w_0_170_s_0_225 = 4.94e-12
+ mcm4l1f_ca_w_0_170_s_0_270 = 3.93e-05  mcm4l1f_cc_w_0_170_s_0_270 = 5.05e-11  mcm4l1f_cf_w_0_170_s_0_270 = 5.74e-12
+ mcm4l1f_ca_w_0_170_s_0_360 = 3.93e-05  mcm4l1f_cc_w_0_170_s_0_360 = 4.20e-11  mcm4l1f_cf_w_0_170_s_0_360 = 7.51e-12
+ mcm4l1f_ca_w_0_170_s_0_450 = 3.93e-05  mcm4l1f_cc_w_0_170_s_0_450 = 3.65e-11  mcm4l1f_cf_w_0_170_s_0_450 = 8.83e-12
+ mcm4l1f_ca_w_0_170_s_0_540 = 3.93e-05  mcm4l1f_cc_w_0_170_s_0_540 = 3.18e-11  mcm4l1f_cf_w_0_170_s_0_540 = 1.05e-11
+ mcm4l1f_ca_w_0_170_s_0_720 = 3.93e-05  mcm4l1f_cc_w_0_170_s_0_720 = 2.55e-11  mcm4l1f_cf_w_0_170_s_0_720 = 1.31e-11
+ mcm4l1f_ca_w_0_170_s_1_080 = 3.93e-05  mcm4l1f_cc_w_0_170_s_1_080 = 1.74e-11  mcm4l1f_cf_w_0_170_s_1_080 = 1.75e-11
+ mcm4l1f_ca_w_0_170_s_1_980 = 3.93e-05  mcm4l1f_cc_w_0_170_s_1_980 = 7.86e-12  mcm4l1f_cf_w_0_170_s_1_980 = 2.44e-11
+ mcm4l1f_ca_w_0_170_s_4_500 = 3.93e-05  mcm4l1f_cc_w_0_170_s_4_500 = 1.21e-12  mcm4l1f_cf_w_0_170_s_4_500 = 3.03e-11
+ mcm4l1f_ca_w_1_360_s_0_180 = 3.93e-05  mcm4l1f_cc_w_1_360_s_0_180 = 8.24e-11  mcm4l1f_cf_w_1_360_s_0_180 = 4.10e-12
+ mcm4l1f_ca_w_1_360_s_0_225 = 3.93e-05  mcm4l1f_cc_w_1_360_s_0_225 = 7.34e-11  mcm4l1f_cf_w_1_360_s_0_225 = 4.94e-12
+ mcm4l1f_ca_w_1_360_s_0_270 = 3.93e-05  mcm4l1f_cc_w_1_360_s_0_270 = 6.63e-11  mcm4l1f_cf_w_1_360_s_0_270 = 5.77e-12
+ mcm4l1f_ca_w_1_360_s_0_360 = 3.93e-05  mcm4l1f_cc_w_1_360_s_0_360 = 5.61e-11  mcm4l1f_cf_w_1_360_s_0_360 = 7.37e-12
+ mcm4l1f_ca_w_1_360_s_0_450 = 3.93e-05  mcm4l1f_cc_w_1_360_s_0_450 = 4.87e-11  mcm4l1f_cf_w_1_360_s_0_450 = 8.93e-12
+ mcm4l1f_ca_w_1_360_s_0_540 = 3.93e-05  mcm4l1f_cc_w_1_360_s_0_540 = 4.31e-11  mcm4l1f_cf_w_1_360_s_0_540 = 1.04e-11
+ mcm4l1f_ca_w_1_360_s_0_720 = 3.93e-05  mcm4l1f_cc_w_1_360_s_0_720 = 3.49e-11  mcm4l1f_cf_w_1_360_s_0_720 = 1.32e-11
+ mcm4l1f_ca_w_1_360_s_1_080 = 3.93e-05  mcm4l1f_cc_w_1_360_s_1_080 = 2.45e-11  mcm4l1f_cf_w_1_360_s_1_080 = 1.81e-11
+ mcm4l1f_ca_w_1_360_s_1_980 = 3.93e-05  mcm4l1f_cc_w_1_360_s_1_980 = 1.16e-11  mcm4l1f_cf_w_1_360_s_1_980 = 2.66e-11
+ mcm4l1f_ca_w_1_360_s_4_500 = 3.93e-05  mcm4l1f_cc_w_1_360_s_4_500 = 1.95e-12  mcm4l1f_cf_w_1_360_s_4_500 = 3.50e-11
+ mcm4l1d_ca_w_0_170_s_0_180 = 5.52e-05  mcm4l1d_cc_w_0_170_s_0_180 = 6.16e-11  mcm4l1d_cf_w_0_170_s_0_180 = 5.72e-12
+ mcm4l1d_ca_w_0_170_s_0_225 = 5.52e-05  mcm4l1d_cc_w_0_170_s_0_225 = 5.36e-11  mcm4l1d_cf_w_0_170_s_0_225 = 6.86e-12
+ mcm4l1d_ca_w_0_170_s_0_270 = 5.52e-05  mcm4l1d_cc_w_0_170_s_0_270 = 4.80e-11  mcm4l1d_cf_w_0_170_s_0_270 = 7.94e-12
+ mcm4l1d_ca_w_0_170_s_0_360 = 5.52e-05  mcm4l1d_cc_w_0_170_s_0_360 = 3.92e-11  mcm4l1d_cf_w_0_170_s_0_360 = 1.03e-11
+ mcm4l1d_ca_w_0_170_s_0_450 = 5.52e-05  mcm4l1d_cc_w_0_170_s_0_450 = 3.35e-11  mcm4l1d_cf_w_0_170_s_0_450 = 1.21e-11
+ mcm4l1d_ca_w_0_170_s_0_540 = 5.52e-05  mcm4l1d_cc_w_0_170_s_0_540 = 2.87e-11  mcm4l1d_cf_w_0_170_s_0_540 = 1.41e-11
+ mcm4l1d_ca_w_0_170_s_0_720 = 5.52e-05  mcm4l1d_cc_w_0_170_s_0_720 = 2.21e-11  mcm4l1d_cf_w_0_170_s_0_720 = 1.74e-11
+ mcm4l1d_ca_w_0_170_s_1_080 = 5.52e-05  mcm4l1d_cc_w_0_170_s_1_080 = 1.41e-11  mcm4l1d_cf_w_0_170_s_1_080 = 2.26e-11
+ mcm4l1d_ca_w_0_170_s_1_980 = 5.52e-05  mcm4l1d_cc_w_0_170_s_1_980 = 5.51e-12  mcm4l1d_cf_w_0_170_s_1_980 = 2.95e-11
+ mcm4l1d_ca_w_0_170_s_4_500 = 5.52e-05  mcm4l1d_cc_w_0_170_s_4_500 = 6.80e-13  mcm4l1d_cf_w_0_170_s_4_500 = 3.40e-11
+ mcm4l1d_ca_w_1_360_s_0_180 = 5.52e-05  mcm4l1d_cc_w_1_360_s_0_180 = 7.79e-11  mcm4l1d_cf_w_1_360_s_0_180 = 5.71e-12
+ mcm4l1d_ca_w_1_360_s_0_225 = 5.52e-05  mcm4l1d_cc_w_1_360_s_0_225 = 6.87e-11  mcm4l1d_cf_w_1_360_s_0_225 = 6.86e-12
+ mcm4l1d_ca_w_1_360_s_0_270 = 5.52e-05  mcm4l1d_cc_w_1_360_s_0_270 = 6.17e-11  mcm4l1d_cf_w_1_360_s_0_270 = 7.98e-12
+ mcm4l1d_ca_w_1_360_s_0_360 = 5.52e-05  mcm4l1d_cc_w_1_360_s_0_360 = 5.14e-11  mcm4l1d_cf_w_1_360_s_0_360 = 1.01e-11
+ mcm4l1d_ca_w_1_360_s_0_450 = 5.52e-05  mcm4l1d_cc_w_1_360_s_0_450 = 4.41e-11  mcm4l1d_cf_w_1_360_s_0_450 = 1.22e-11
+ mcm4l1d_ca_w_1_360_s_0_540 = 5.52e-05  mcm4l1d_cc_w_1_360_s_0_540 = 3.85e-11  mcm4l1d_cf_w_1_360_s_0_540 = 1.42e-11
+ mcm4l1d_ca_w_1_360_s_0_720 = 5.52e-05  mcm4l1d_cc_w_1_360_s_0_720 = 3.04e-11  mcm4l1d_cf_w_1_360_s_0_720 = 1.77e-11
+ mcm4l1d_ca_w_1_360_s_1_080 = 5.52e-05  mcm4l1d_cc_w_1_360_s_1_080 = 2.03e-11  mcm4l1d_cf_w_1_360_s_1_080 = 2.35e-11
+ mcm4l1d_ca_w_1_360_s_1_980 = 5.52e-05  mcm4l1d_cc_w_1_360_s_1_980 = 8.67e-12  mcm4l1d_cf_w_1_360_s_1_980 = 3.23e-11
+ mcm4l1d_ca_w_1_360_s_4_500 = 5.52e-05  mcm4l1d_cc_w_1_360_s_4_500 = 1.23e-12  mcm4l1d_cf_w_1_360_s_4_500 = 3.92e-11
+ mcm4l1p1_ca_w_0_170_s_0_180 = 7.44e-05  mcm4l1p1_cc_w_0_170_s_0_180 = 5.92e-11  mcm4l1p1_cf_w_0_170_s_0_180 = 7.63e-12
+ mcm4l1p1_ca_w_0_170_s_0_225 = 7.44e-05  mcm4l1p1_cc_w_0_170_s_0_225 = 5.11e-11  mcm4l1p1_cf_w_0_170_s_0_225 = 9.11e-12
+ mcm4l1p1_ca_w_0_170_s_0_270 = 7.44e-05  mcm4l1p1_cc_w_0_170_s_0_270 = 4.53e-11  mcm4l1p1_cf_w_0_170_s_0_270 = 1.05e-11
+ mcm4l1p1_ca_w_0_170_s_0_360 = 7.44e-05  mcm4l1p1_cc_w_0_170_s_0_360 = 3.63e-11  mcm4l1p1_cf_w_0_170_s_0_360 = 1.35e-11
+ mcm4l1p1_ca_w_0_170_s_0_450 = 7.44e-05  mcm4l1p1_cc_w_0_170_s_0_450 = 3.06e-11  mcm4l1p1_cf_w_0_170_s_0_450 = 1.57e-11
+ mcm4l1p1_ca_w_0_170_s_0_540 = 7.44e-05  mcm4l1p1_cc_w_0_170_s_0_540 = 2.56e-11  mcm4l1p1_cf_w_0_170_s_0_540 = 1.82e-11
+ mcm4l1p1_ca_w_0_170_s_0_720 = 7.44e-05  mcm4l1p1_cc_w_0_170_s_0_720 = 1.90e-11  mcm4l1p1_cf_w_0_170_s_0_720 = 2.21e-11
+ mcm4l1p1_ca_w_0_170_s_1_080 = 7.44e-05  mcm4l1p1_cc_w_0_170_s_1_080 = 1.14e-11  mcm4l1p1_cf_w_0_170_s_1_080 = 2.76e-11
+ mcm4l1p1_ca_w_0_170_s_1_980 = 7.44e-05  mcm4l1p1_cc_w_0_170_s_1_980 = 3.96e-12  mcm4l1p1_cf_w_0_170_s_1_980 = 3.41e-11
+ mcm4l1p1_ca_w_0_170_s_4_500 = 7.44e-05  mcm4l1p1_cc_w_0_170_s_4_500 = 4.30e-13  mcm4l1p1_cf_w_0_170_s_4_500 = 3.74e-11
+ mcm4l1p1_ca_w_1_360_s_0_180 = 7.44e-05  mcm4l1p1_cc_w_1_360_s_0_180 = 7.40e-11  mcm4l1p1_cf_w_1_360_s_0_180 = 7.67e-12
+ mcm4l1p1_ca_w_1_360_s_0_225 = 7.44e-05  mcm4l1p1_cc_w_1_360_s_0_225 = 6.48e-11  mcm4l1p1_cf_w_1_360_s_0_225 = 9.17e-12
+ mcm4l1p1_ca_w_1_360_s_0_270 = 7.44e-05  mcm4l1p1_cc_w_1_360_s_0_270 = 5.78e-11  mcm4l1p1_cf_w_1_360_s_0_270 = 1.06e-11
+ mcm4l1p1_ca_w_1_360_s_0_360 = 7.44e-05  mcm4l1p1_cc_w_1_360_s_0_360 = 4.76e-11  mcm4l1p1_cf_w_1_360_s_0_360 = 1.34e-11
+ mcm4l1p1_ca_w_1_360_s_0_450 = 7.44e-05  mcm4l1p1_cc_w_1_360_s_0_450 = 4.03e-11  mcm4l1p1_cf_w_1_360_s_0_450 = 1.60e-11
+ mcm4l1p1_ca_w_1_360_s_0_540 = 7.44e-05  mcm4l1p1_cc_w_1_360_s_0_540 = 3.48e-11  mcm4l1p1_cf_w_1_360_s_0_540 = 1.83e-11
+ mcm4l1p1_ca_w_1_360_s_0_720 = 7.44e-05  mcm4l1p1_cc_w_1_360_s_0_720 = 2.68e-11  mcm4l1p1_cf_w_1_360_s_0_720 = 2.25e-11
+ mcm4l1p1_ca_w_1_360_s_1_080 = 7.44e-05  mcm4l1p1_cc_w_1_360_s_1_080 = 1.72e-11  mcm4l1p1_cf_w_1_360_s_1_080 = 2.89e-11
+ mcm4l1p1_ca_w_1_360_s_1_980 = 7.44e-05  mcm4l1p1_cc_w_1_360_s_1_980 = 6.80e-12  mcm4l1p1_cf_w_1_360_s_1_980 = 3.75e-11
+ mcm4l1p1_ca_w_1_360_s_4_500 = 7.44e-05  mcm4l1p1_cc_w_1_360_s_4_500 = 8.25e-13  mcm4l1p1_cf_w_1_360_s_4_500 = 4.32e-11
+ mcm5l1f_ca_w_0_170_s_0_180 = 3.63e-05  mcm5l1f_cc_w_0_170_s_0_180 = 6.42e-11  mcm5l1f_cf_w_0_170_s_0_180 = 3.81e-12
+ mcm5l1f_ca_w_0_170_s_0_225 = 3.63e-05  mcm5l1f_cc_w_0_170_s_0_225 = 5.63e-11  mcm5l1f_cf_w_0_170_s_0_225 = 4.58e-12
+ mcm5l1f_ca_w_0_170_s_0_270 = 3.63e-05  mcm5l1f_cc_w_0_170_s_0_270 = 5.11e-11  mcm5l1f_cf_w_0_170_s_0_270 = 5.31e-12
+ mcm5l1f_ca_w_0_170_s_0_360 = 3.63e-05  mcm5l1f_cc_w_0_170_s_0_360 = 4.26e-11  mcm5l1f_cf_w_0_170_s_0_360 = 6.97e-12
+ mcm5l1f_ca_w_0_170_s_0_450 = 3.63e-05  mcm5l1f_cc_w_0_170_s_0_450 = 3.72e-11  mcm5l1f_cf_w_0_170_s_0_450 = 8.20e-12
+ mcm5l1f_ca_w_0_170_s_0_540 = 3.63e-05  mcm5l1f_cc_w_0_170_s_0_540 = 3.26e-11  mcm5l1f_cf_w_0_170_s_0_540 = 9.75e-12
+ mcm5l1f_ca_w_0_170_s_0_720 = 3.63e-05  mcm5l1f_cc_w_0_170_s_0_720 = 2.63e-11  mcm5l1f_cf_w_0_170_s_0_720 = 1.23e-11
+ mcm5l1f_ca_w_0_170_s_1_080 = 3.63e-05  mcm5l1f_cc_w_0_170_s_1_080 = 1.84e-11  mcm5l1f_cf_w_0_170_s_1_080 = 1.65e-11
+ mcm5l1f_ca_w_0_170_s_1_980 = 3.63e-05  mcm5l1f_cc_w_0_170_s_1_980 = 8.93e-12  mcm5l1f_cf_w_0_170_s_1_980 = 2.32e-11
+ mcm5l1f_ca_w_0_170_s_4_500 = 3.63e-05  mcm5l1f_cc_w_0_170_s_4_500 = 1.73e-12  mcm5l1f_cf_w_0_170_s_4_500 = 2.95e-11
+ mcm5l1f_ca_w_1_360_s_0_180 = 3.63e-05  mcm5l1f_cc_w_1_360_s_0_180 = 8.44e-11  mcm5l1f_cf_w_1_360_s_0_180 = 3.80e-12
+ mcm5l1f_ca_w_1_360_s_0_225 = 3.63e-05  mcm5l1f_cc_w_1_360_s_0_225 = 7.52e-11  mcm5l1f_cf_w_1_360_s_0_225 = 4.58e-12
+ mcm5l1f_ca_w_1_360_s_0_270 = 3.63e-05  mcm5l1f_cc_w_1_360_s_0_270 = 6.81e-11  mcm5l1f_cf_w_1_360_s_0_270 = 5.34e-12
+ mcm5l1f_ca_w_1_360_s_0_360 = 3.63e-05  mcm5l1f_cc_w_1_360_s_0_360 = 5.80e-11  mcm5l1f_cf_w_1_360_s_0_360 = 6.83e-12
+ mcm5l1f_ca_w_1_360_s_0_450 = 3.63e-05  mcm5l1f_cc_w_1_360_s_0_450 = 5.07e-11  mcm5l1f_cf_w_1_360_s_0_450 = 8.29e-12
+ mcm5l1f_ca_w_1_360_s_0_540 = 3.63e-05  mcm5l1f_cc_w_1_360_s_0_540 = 4.52e-11  mcm5l1f_cf_w_1_360_s_0_540 = 9.69e-12
+ mcm5l1f_ca_w_1_360_s_0_720 = 3.63e-05  mcm5l1f_cc_w_1_360_s_0_720 = 3.71e-11  mcm5l1f_cf_w_1_360_s_0_720 = 1.23e-11
+ mcm5l1f_ca_w_1_360_s_1_080 = 3.63e-05  mcm5l1f_cc_w_1_360_s_1_080 = 2.67e-11  mcm5l1f_cf_w_1_360_s_1_080 = 1.69e-11
+ mcm5l1f_ca_w_1_360_s_1_980 = 3.63e-05  mcm5l1f_cc_w_1_360_s_1_980 = 1.37e-11  mcm5l1f_cf_w_1_360_s_1_980 = 2.52e-11
+ mcm5l1f_ca_w_1_360_s_4_500 = 3.63e-05  mcm5l1f_cc_w_1_360_s_4_500 = 3.01e-12  mcm5l1f_cf_w_1_360_s_4_500 = 3.44e-11
+ mcm5l1d_ca_w_0_170_s_0_180 = 5.22e-05  mcm5l1d_cc_w_0_170_s_0_180 = 6.19e-11  mcm5l1d_cf_w_0_170_s_0_180 = 5.42e-12
+ mcm5l1d_ca_w_0_170_s_0_225 = 5.22e-05  mcm5l1d_cc_w_0_170_s_0_225 = 5.40e-11  mcm5l1d_cf_w_0_170_s_0_225 = 6.50e-12
+ mcm5l1d_ca_w_0_170_s_0_270 = 5.22e-05  mcm5l1d_cc_w_0_170_s_0_270 = 4.85e-11  mcm5l1d_cf_w_0_170_s_0_270 = 7.53e-12
+ mcm5l1d_ca_w_0_170_s_0_360 = 5.22e-05  mcm5l1d_cc_w_0_170_s_0_360 = 3.98e-11  mcm5l1d_cf_w_0_170_s_0_360 = 9.76e-12
+ mcm5l1d_ca_w_0_170_s_0_450 = 5.22e-05  mcm5l1d_cc_w_0_170_s_0_450 = 3.42e-11  mcm5l1d_cf_w_0_170_s_0_450 = 1.15e-11
+ mcm5l1d_ca_w_0_170_s_0_540 = 5.22e-05  mcm5l1d_cc_w_0_170_s_0_540 = 2.94e-11  mcm5l1d_cf_w_0_170_s_0_540 = 1.34e-11
+ mcm5l1d_ca_w_0_170_s_0_720 = 5.22e-05  mcm5l1d_cc_w_0_170_s_0_720 = 2.29e-11  mcm5l1d_cf_w_0_170_s_0_720 = 1.67e-11
+ mcm5l1d_ca_w_0_170_s_1_080 = 5.22e-05  mcm5l1d_cc_w_0_170_s_1_080 = 1.50e-11  mcm5l1d_cf_w_0_170_s_1_080 = 2.17e-11
+ mcm5l1d_ca_w_0_170_s_1_980 = 5.22e-05  mcm5l1d_cc_w_0_170_s_1_980 = 6.34e-12  mcm5l1d_cf_w_0_170_s_1_980 = 2.86e-11
+ mcm5l1d_ca_w_0_170_s_4_500 = 5.22e-05  mcm5l1d_cc_w_0_170_s_4_500 = 1.02e-12  mcm5l1d_cf_w_0_170_s_4_500 = 3.35e-11
+ mcm5l1d_ca_w_1_360_s_0_180 = 5.22e-05  mcm5l1d_cc_w_1_360_s_0_180 = 7.96e-11  mcm5l1d_cf_w_1_360_s_0_180 = 5.41e-12
+ mcm5l1d_ca_w_1_360_s_0_225 = 5.22e-05  mcm5l1d_cc_w_1_360_s_0_225 = 7.06e-11  mcm5l1d_cf_w_1_360_s_0_225 = 6.50e-12
+ mcm5l1d_ca_w_1_360_s_0_270 = 5.22e-05  mcm5l1d_cc_w_1_360_s_0_270 = 6.36e-11  mcm5l1d_cf_w_1_360_s_0_270 = 7.57e-12
+ mcm5l1d_ca_w_1_360_s_0_360 = 5.22e-05  mcm5l1d_cc_w_1_360_s_0_360 = 5.34e-11  mcm5l1d_cf_w_1_360_s_0_360 = 9.62e-12
+ mcm5l1d_ca_w_1_360_s_0_450 = 5.22e-05  mcm5l1d_cc_w_1_360_s_0_450 = 4.61e-11  mcm5l1d_cf_w_1_360_s_0_450 = 1.16e-11
+ mcm5l1d_ca_w_1_360_s_0_540 = 5.22e-05  mcm5l1d_cc_w_1_360_s_0_540 = 4.06e-11  mcm5l1d_cf_w_1_360_s_0_540 = 1.34e-11
+ mcm5l1d_ca_w_1_360_s_0_720 = 5.22e-05  mcm5l1d_cc_w_1_360_s_0_720 = 3.25e-11  mcm5l1d_cf_w_1_360_s_0_720 = 1.68e-11
+ mcm5l1d_ca_w_1_360_s_1_080 = 5.22e-05  mcm5l1d_cc_w_1_360_s_1_080 = 2.24e-11  mcm5l1d_cf_w_1_360_s_1_080 = 2.25e-11
+ mcm5l1d_ca_w_1_360_s_1_980 = 5.22e-05  mcm5l1d_cc_w_1_360_s_1_980 = 1.04e-11  mcm5l1d_cf_w_1_360_s_1_980 = 3.14e-11
+ mcm5l1d_ca_w_1_360_s_4_500 = 5.22e-05  mcm5l1d_cc_w_1_360_s_4_500 = 1.99e-12  mcm5l1d_cf_w_1_360_s_4_500 = 3.91e-11
+ mcm5l1p1_ca_w_0_170_s_0_180 = 7.15e-05  mcm5l1p1_cc_w_0_170_s_0_180 = 5.95e-11  mcm5l1p1_cf_w_0_170_s_0_180 = 7.33e-12
+ mcm5l1p1_ca_w_0_170_s_0_225 = 7.15e-05  mcm5l1p1_cc_w_0_170_s_0_225 = 5.15e-11  mcm5l1p1_cf_w_0_170_s_0_225 = 8.74e-12
+ mcm5l1p1_ca_w_0_170_s_0_270 = 7.15e-05  mcm5l1p1_cc_w_0_170_s_0_270 = 4.58e-11  mcm5l1p1_cf_w_0_170_s_0_270 = 1.01e-11
+ mcm5l1p1_ca_w_0_170_s_0_360 = 7.15e-05  mcm5l1p1_cc_w_0_170_s_0_360 = 3.69e-11  mcm5l1p1_cf_w_0_170_s_0_360 = 1.30e-11
+ mcm5l1p1_ca_w_0_170_s_0_450 = 7.15e-05  mcm5l1p1_cc_w_0_170_s_0_450 = 3.12e-11  mcm5l1p1_cf_w_0_170_s_0_450 = 1.51e-11
+ mcm5l1p1_ca_w_0_170_s_0_540 = 7.15e-05  mcm5l1p1_cc_w_0_170_s_0_540 = 2.63e-11  mcm5l1p1_cf_w_0_170_s_0_540 = 1.76e-11
+ mcm5l1p1_ca_w_0_170_s_0_720 = 7.15e-05  mcm5l1p1_cc_w_0_170_s_0_720 = 1.98e-11  mcm5l1p1_cf_w_0_170_s_0_720 = 2.14e-11
+ mcm5l1p1_ca_w_0_170_s_1_080 = 7.15e-05  mcm5l1p1_cc_w_0_170_s_1_080 = 1.21e-11  mcm5l1p1_cf_w_0_170_s_1_080 = 2.69e-11
+ mcm5l1p1_ca_w_0_170_s_1_980 = 7.15e-05  mcm5l1p1_cc_w_0_170_s_1_980 = 4.60e-12  mcm5l1p1_cf_w_0_170_s_1_980 = 3.34e-11
+ mcm5l1p1_ca_w_0_170_s_4_500 = 7.15e-05  mcm5l1p1_cc_w_0_170_s_4_500 = 6.63e-13  mcm5l1p1_cf_w_0_170_s_4_500 = 3.71e-11
+ mcm5l1p1_ca_w_1_360_s_0_180 = 7.15e-05  mcm5l1p1_cc_w_1_360_s_0_180 = 7.58e-11  mcm5l1p1_cf_w_1_360_s_0_180 = 7.37e-12
+ mcm5l1p1_ca_w_1_360_s_0_225 = 7.15e-05  mcm5l1p1_cc_w_1_360_s_0_225 = 6.66e-11  mcm5l1p1_cf_w_1_360_s_0_225 = 8.81e-12
+ mcm5l1p1_ca_w_1_360_s_0_270 = 7.15e-05  mcm5l1p1_cc_w_1_360_s_0_270 = 5.96e-11  mcm5l1p1_cf_w_1_360_s_0_270 = 1.02e-11
+ mcm5l1p1_ca_w_1_360_s_0_360 = 7.15e-05  mcm5l1p1_cc_w_1_360_s_0_360 = 4.95e-11  mcm5l1p1_cf_w_1_360_s_0_360 = 1.29e-11
+ mcm5l1p1_ca_w_1_360_s_0_450 = 7.15e-05  mcm5l1p1_cc_w_1_360_s_0_450 = 4.23e-11  mcm5l1p1_cf_w_1_360_s_0_450 = 1.54e-11
+ mcm5l1p1_ca_w_1_360_s_0_540 = 7.15e-05  mcm5l1p1_cc_w_1_360_s_0_540 = 3.68e-11  mcm5l1p1_cf_w_1_360_s_0_540 = 1.77e-11
+ mcm5l1p1_ca_w_1_360_s_0_720 = 7.15e-05  mcm5l1p1_cc_w_1_360_s_0_720 = 2.89e-11  mcm5l1p1_cf_w_1_360_s_0_720 = 2.18e-11
+ mcm5l1p1_ca_w_1_360_s_1_080 = 7.15e-05  mcm5l1p1_cc_w_1_360_s_1_080 = 1.92e-11  mcm5l1p1_cf_w_1_360_s_1_080 = 2.81e-11
+ mcm5l1p1_ca_w_1_360_s_1_980 = 7.15e-05  mcm5l1p1_cc_w_1_360_s_1_980 = 8.41e-12  mcm5l1p1_cf_w_1_360_s_1_980 = 3.69e-11
+ mcm5l1p1_ca_w_1_360_s_4_500 = 7.15e-05  mcm5l1p1_cc_w_1_360_s_4_500 = 1.47e-12  mcm5l1p1_cf_w_1_360_s_4_500 = 4.34e-11
+ mcrdll1f_ca_w_0_170_s_0_180 = 3.17e-05  mcrdll1f_cc_w_0_170_s_0_180 = 6.47e-11  mcrdll1f_cf_w_0_170_s_0_180 = 3.32e-12
+ mcrdll1f_ca_w_0_170_s_0_225 = 3.17e-05  mcrdll1f_cc_w_0_170_s_0_225 = 5.70e-11  mcrdll1f_cf_w_0_170_s_0_225 = 3.99e-12
+ mcrdll1f_ca_w_0_170_s_0_270 = 3.17e-05  mcrdll1f_cc_w_0_170_s_0_270 = 5.18e-11  mcrdll1f_cf_w_0_170_s_0_270 = 4.65e-12
+ mcrdll1f_ca_w_0_170_s_0_360 = 3.17e-05  mcrdll1f_cc_w_0_170_s_0_360 = 4.34e-11  mcrdll1f_cf_w_0_170_s_0_360 = 6.10e-12
+ mcrdll1f_ca_w_0_170_s_0_450 = 3.17e-05  mcrdll1f_cc_w_0_170_s_0_450 = 3.84e-11  mcrdll1f_cf_w_0_170_s_0_450 = 7.18e-12
+ mcrdll1f_ca_w_0_170_s_0_540 = 3.17e-05  mcrdll1f_cc_w_0_170_s_0_540 = 3.38e-11  mcrdll1f_cf_w_0_170_s_0_540 = 8.59e-12
+ mcrdll1f_ca_w_0_170_s_0_720 = 3.17e-05  mcrdll1f_cc_w_0_170_s_0_720 = 2.77e-11  mcrdll1f_cf_w_0_170_s_0_720 = 1.09e-11
+ mcrdll1f_ca_w_0_170_s_1_080 = 3.17e-05  mcrdll1f_cc_w_0_170_s_1_080 = 2.00e-11  mcrdll1f_cf_w_0_170_s_1_080 = 1.48e-11
+ mcrdll1f_ca_w_0_170_s_1_980 = 3.17e-05  mcrdll1f_cc_w_0_170_s_1_980 = 1.09e-11  mcrdll1f_cf_w_0_170_s_1_980 = 2.11e-11
+ mcrdll1f_ca_w_0_170_s_4_500 = 3.17e-05  mcrdll1f_cc_w_0_170_s_4_500 = 3.01e-12  mcrdll1f_cf_w_0_170_s_4_500 = 2.80e-11
+ mcrdll1f_ca_w_1_360_s_0_180 = 3.17e-05  mcrdll1f_cc_w_1_360_s_0_180 = 8.73e-11  mcrdll1f_cf_w_1_360_s_0_180 = 3.32e-12
+ mcrdll1f_ca_w_1_360_s_0_225 = 3.17e-05  mcrdll1f_cc_w_1_360_s_0_225 = 7.82e-11  mcrdll1f_cf_w_1_360_s_0_225 = 4.00e-12
+ mcrdll1f_ca_w_1_360_s_0_270 = 3.17e-05  mcrdll1f_cc_w_1_360_s_0_270 = 7.14e-11  mcrdll1f_cf_w_1_360_s_0_270 = 4.67e-12
+ mcrdll1f_ca_w_1_360_s_0_360 = 3.17e-05  mcrdll1f_cc_w_1_360_s_0_360 = 6.13e-11  mcrdll1f_cf_w_1_360_s_0_360 = 5.98e-12
+ mcrdll1f_ca_w_1_360_s_0_450 = 3.17e-05  mcrdll1f_cc_w_1_360_s_0_450 = 5.42e-11  mcrdll1f_cf_w_1_360_s_0_450 = 7.26e-12
+ mcrdll1f_ca_w_1_360_s_0_540 = 3.17e-05  mcrdll1f_cc_w_1_360_s_0_540 = 4.87e-11  mcrdll1f_cf_w_1_360_s_0_540 = 8.50e-12
+ mcrdll1f_ca_w_1_360_s_0_720 = 3.17e-05  mcrdll1f_cc_w_1_360_s_0_720 = 4.07e-11  mcrdll1f_cf_w_1_360_s_0_720 = 1.08e-11
+ mcrdll1f_ca_w_1_360_s_1_080 = 3.17e-05  mcrdll1f_cc_w_1_360_s_1_080 = 3.07e-11  mcrdll1f_cf_w_1_360_s_1_080 = 1.50e-11
+ mcrdll1f_ca_w_1_360_s_1_980 = 3.17e-05  mcrdll1f_cc_w_1_360_s_1_980 = 1.78e-11  mcrdll1f_cf_w_1_360_s_1_980 = 2.29e-11
+ mcrdll1f_ca_w_1_360_s_4_500 = 3.17e-05  mcrdll1f_cc_w_1_360_s_4_500 = 5.84e-12  mcrdll1f_cf_w_1_360_s_4_500 = 3.29e-11
+ mcrdll1d_ca_w_0_170_s_0_180 = 4.76e-05  mcrdll1d_cc_w_0_170_s_0_180 = 6.25e-11  mcrdll1d_cf_w_0_170_s_0_180 = 4.94e-12
+ mcrdll1d_ca_w_0_170_s_0_225 = 4.76e-05  mcrdll1d_cc_w_0_170_s_0_225 = 5.47e-11  mcrdll1d_cf_w_0_170_s_0_225 = 5.92e-12
+ mcrdll1d_ca_w_0_170_s_0_270 = 4.76e-05  mcrdll1d_cc_w_0_170_s_0_270 = 4.93e-11  mcrdll1d_cf_w_0_170_s_0_270 = 6.88e-12
+ mcrdll1d_ca_w_0_170_s_0_360 = 4.76e-05  mcrdll1d_cc_w_0_170_s_0_360 = 4.07e-11  mcrdll1d_cf_w_0_170_s_0_360 = 8.93e-12
+ mcrdll1d_ca_w_0_170_s_0_450 = 4.76e-05  mcrdll1d_cc_w_0_170_s_0_450 = 3.53e-11  mcrdll1d_cf_w_0_170_s_0_450 = 1.05e-11
+ mcrdll1d_ca_w_0_170_s_0_540 = 4.76e-05  mcrdll1d_cc_w_0_170_s_0_540 = 3.05e-11  mcrdll1d_cf_w_0_170_s_0_540 = 1.24e-11
+ mcrdll1d_ca_w_0_170_s_0_720 = 4.76e-05  mcrdll1d_cc_w_0_170_s_0_720 = 2.42e-11  mcrdll1d_cf_w_0_170_s_0_720 = 1.54e-11
+ mcrdll1d_ca_w_0_170_s_1_080 = 4.76e-05  mcrdll1d_cc_w_0_170_s_1_080 = 1.64e-11  mcrdll1d_cf_w_0_170_s_1_080 = 2.03e-11
+ mcrdll1d_ca_w_0_170_s_1_980 = 4.76e-05  mcrdll1d_cc_w_0_170_s_1_980 = 7.85e-12  mcrdll1d_cf_w_0_170_s_1_980 = 2.71e-11
+ mcrdll1d_ca_w_0_170_s_4_500 = 4.76e-05  mcrdll1d_cc_w_0_170_s_4_500 = 1.86e-12  mcrdll1d_cf_w_0_170_s_4_500 = 3.26e-11
+ mcrdll1d_ca_w_1_360_s_0_180 = 4.76e-05  mcrdll1d_cc_w_1_360_s_0_180 = 8.26e-11  mcrdll1d_cf_w_1_360_s_0_180 = 4.93e-12
+ mcrdll1d_ca_w_1_360_s_0_225 = 4.76e-05  mcrdll1d_cc_w_1_360_s_0_225 = 7.36e-11  mcrdll1d_cf_w_1_360_s_0_225 = 5.92e-12
+ mcrdll1d_ca_w_1_360_s_0_270 = 4.76e-05  mcrdll1d_cc_w_1_360_s_0_270 = 6.67e-11  mcrdll1d_cf_w_1_360_s_0_270 = 6.90e-12
+ mcrdll1d_ca_w_1_360_s_0_360 = 4.76e-05  mcrdll1d_cc_w_1_360_s_0_360 = 5.66e-11  mcrdll1d_cf_w_1_360_s_0_360 = 8.80e-12
+ mcrdll1d_ca_w_1_360_s_0_450 = 4.76e-05  mcrdll1d_cc_w_1_360_s_0_450 = 4.95e-11  mcrdll1d_cf_w_1_360_s_0_450 = 1.06e-11
+ mcrdll1d_ca_w_1_360_s_0_540 = 4.76e-05  mcrdll1d_cc_w_1_360_s_0_540 = 4.40e-11  mcrdll1d_cf_w_1_360_s_0_540 = 1.23e-11
+ mcrdll1d_ca_w_1_360_s_0_720 = 4.76e-05  mcrdll1d_cc_w_1_360_s_0_720 = 3.61e-11  mcrdll1d_cf_w_1_360_s_0_720 = 1.55e-11
+ mcrdll1d_ca_w_1_360_s_1_080 = 4.76e-05  mcrdll1d_cc_w_1_360_s_1_080 = 2.62e-11  mcrdll1d_cf_w_1_360_s_1_080 = 2.08e-11
+ mcrdll1d_ca_w_1_360_s_1_980 = 4.76e-05  mcrdll1d_cc_w_1_360_s_1_980 = 1.41e-11  mcrdll1d_cf_w_1_360_s_1_980 = 2.97e-11
+ mcrdll1d_ca_w_1_360_s_4_500 = 4.76e-05  mcrdll1d_cc_w_1_360_s_4_500 = 4.20e-12  mcrdll1d_cf_w_1_360_s_4_500 = 3.86e-11
+ mcrdll1p1_ca_w_0_170_s_0_180 = 6.68e-05  mcrdll1p1_cc_w_0_170_s_0_180 = 6.01e-11  mcrdll1p1_cf_w_0_170_s_0_180 = 6.85e-12
+ mcrdll1p1_ca_w_0_170_s_0_225 = 6.68e-05  mcrdll1p1_cc_w_0_170_s_0_225 = 5.22e-11  mcrdll1p1_cf_w_0_170_s_0_225 = 8.17e-12
+ mcrdll1p1_ca_w_0_170_s_0_270 = 6.68e-05  mcrdll1p1_cc_w_0_170_s_0_270 = 4.66e-11  mcrdll1p1_cf_w_0_170_s_0_270 = 9.47e-12
+ mcrdll1p1_ca_w_0_170_s_0_360 = 6.68e-05  mcrdll1p1_cc_w_0_170_s_0_360 = 3.77e-11  mcrdll1p1_cf_w_0_170_s_0_360 = 1.21e-11
+ mcrdll1p1_ca_w_0_170_s_0_450 = 6.68e-05  mcrdll1p1_cc_w_0_170_s_0_450 = 3.22e-11  mcrdll1p1_cf_w_0_170_s_0_450 = 1.42e-11
+ mcrdll1p1_ca_w_0_170_s_0_540 = 6.68e-05  mcrdll1p1_cc_w_0_170_s_0_540 = 2.73e-11  mcrdll1p1_cf_w_0_170_s_0_540 = 1.66e-11
+ mcrdll1p1_ca_w_0_170_s_0_720 = 6.68e-05  mcrdll1p1_cc_w_0_170_s_0_720 = 2.09e-11  mcrdll1p1_cf_w_0_170_s_0_720 = 2.03e-11
+ mcrdll1p1_ca_w_0_170_s_1_080 = 6.68e-05  mcrdll1p1_cc_w_0_170_s_1_080 = 1.33e-11  mcrdll1p1_cf_w_0_170_s_1_080 = 2.57e-11
+ mcrdll1p1_ca_w_0_170_s_1_980 = 6.68e-05  mcrdll1p1_cc_w_0_170_s_1_980 = 5.79e-12  mcrdll1p1_cf_w_0_170_s_1_980 = 3.23e-11
+ mcrdll1p1_ca_w_0_170_s_4_500 = 6.68e-05  mcrdll1p1_cc_w_0_170_s_4_500 = 1.26e-12  mcrdll1p1_cf_w_0_170_s_4_500 = 3.66e-11
+ mcrdll1p1_ca_w_1_360_s_0_180 = 6.68e-05  mcrdll1p1_cc_w_1_360_s_0_180 = 7.87e-11  mcrdll1p1_cf_w_1_360_s_0_180 = 6.91e-12
+ mcrdll1p1_ca_w_1_360_s_0_225 = 6.68e-05  mcrdll1p1_cc_w_1_360_s_0_225 = 6.98e-11  mcrdll1p1_cf_w_1_360_s_0_225 = 8.26e-12
+ mcrdll1p1_ca_w_1_360_s_0_270 = 6.68e-05  mcrdll1p1_cc_w_1_360_s_0_270 = 6.28e-11  mcrdll1p1_cf_w_1_360_s_0_270 = 9.57e-12
+ mcrdll1p1_ca_w_1_360_s_0_360 = 6.68e-05  mcrdll1p1_cc_w_1_360_s_0_360 = 5.27e-11  mcrdll1p1_cf_w_1_360_s_0_360 = 1.21e-11
+ mcrdll1p1_ca_w_1_360_s_0_450 = 6.68e-05  mcrdll1p1_cc_w_1_360_s_0_450 = 4.56e-11  mcrdll1p1_cf_w_1_360_s_0_450 = 1.44e-11
+ mcrdll1p1_ca_w_1_360_s_0_540 = 6.68e-05  mcrdll1p1_cc_w_1_360_s_0_540 = 4.02e-11  mcrdll1p1_cf_w_1_360_s_0_540 = 1.66e-11
+ mcrdll1p1_ca_w_1_360_s_0_720 = 6.68e-05  mcrdll1p1_cc_w_1_360_s_0_720 = 3.24e-11  mcrdll1p1_cf_w_1_360_s_0_720 = 2.05e-11
+ mcrdll1p1_ca_w_1_360_s_1_080 = 6.68e-05  mcrdll1p1_cc_w_1_360_s_1_080 = 2.28e-11  mcrdll1p1_cf_w_1_360_s_1_080 = 2.67e-11
+ mcrdll1p1_ca_w_1_360_s_1_980 = 6.68e-05  mcrdll1p1_cc_w_1_360_s_1_980 = 1.16e-11  mcrdll1p1_cf_w_1_360_s_1_980 = 3.58e-11
+ mcrdll1p1_ca_w_1_360_s_4_500 = 6.68e-05  mcrdll1p1_cc_w_1_360_s_4_500 = 3.25e-12  mcrdll1p1_cf_w_1_360_s_4_500 = 4.36e-11
+ mcm2m1f_ca_w_0_140_s_0_140 = 1.01e-04  mcm2m1f_cc_w_0_140_s_0_140 = 7.97e-11  mcm2m1f_cf_w_0_140_s_0_140 = 7.94e-12
+ mcm2m1f_ca_w_0_140_s_0_175 = 1.01e-04  mcm2m1f_cc_w_0_140_s_0_175 = 7.82e-11  mcm2m1f_cf_w_0_140_s_0_175 = 9.49e-12
+ mcm2m1f_ca_w_0_140_s_0_210 = 1.01e-04  mcm2m1f_cc_w_0_140_s_0_210 = 7.42e-11  mcm2m1f_cf_w_0_140_s_0_210 = 1.11e-11
+ mcm2m1f_ca_w_0_140_s_0_280 = 1.01e-04  mcm2m1f_cc_w_0_140_s_0_280 = 6.48e-11  mcm2m1f_cf_w_0_140_s_0_280 = 1.40e-11
+ mcm2m1f_ca_w_0_140_s_0_350 = 1.01e-04  mcm2m1f_cc_w_0_140_s_0_350 = 5.51e-11  mcm2m1f_cf_w_0_140_s_0_350 = 1.68e-11
+ mcm2m1f_ca_w_0_140_s_0_420 = 1.01e-04  mcm2m1f_cc_w_0_140_s_0_420 = 4.68e-11  mcm2m1f_cf_w_0_140_s_0_420 = 1.96e-11
+ mcm2m1f_ca_w_0_140_s_0_560 = 1.01e-04  mcm2m1f_cc_w_0_140_s_0_560 = 3.51e-11  mcm2m1f_cf_w_0_140_s_0_560 = 2.43e-11
+ mcm2m1f_ca_w_0_140_s_0_840 = 1.01e-04  mcm2m1f_cc_w_0_140_s_0_840 = 2.15e-11  mcm2m1f_cf_w_0_140_s_0_840 = 3.20e-11
+ mcm2m1f_ca_w_0_140_s_1_540 = 1.01e-04  mcm2m1f_cc_w_0_140_s_1_540 = 7.57e-12  mcm2m1f_cf_w_0_140_s_1_540 = 4.28e-11
+ mcm2m1f_ca_w_0_140_s_3_500 = 1.01e-04  mcm2m1f_cc_w_0_140_s_3_500 = 6.70e-13  mcm2m1f_cf_w_0_140_s_3_500 = 4.94e-11
+ mcm2m1f_ca_w_1_120_s_0_140 = 1.01e-04  mcm2m1f_cc_w_1_120_s_0_140 = 9.21e-11  mcm2m1f_cf_w_1_120_s_0_140 = 8.00e-12
+ mcm2m1f_ca_w_1_120_s_0_175 = 1.01e-04  mcm2m1f_cc_w_1_120_s_0_175 = 8.90e-11  mcm2m1f_cf_w_1_120_s_0_175 = 9.57e-12
+ mcm2m1f_ca_w_1_120_s_0_210 = 1.01e-04  mcm2m1f_cc_w_1_120_s_0_210 = 8.41e-11  mcm2m1f_cf_w_1_120_s_0_210 = 1.11e-11
+ mcm2m1f_ca_w_1_120_s_0_280 = 1.01e-04  mcm2m1f_cc_w_1_120_s_0_280 = 7.32e-11  mcm2m1f_cf_w_1_120_s_0_280 = 1.41e-11
+ mcm2m1f_ca_w_1_120_s_0_350 = 1.01e-04  mcm2m1f_cc_w_1_120_s_0_350 = 6.23e-11  mcm2m1f_cf_w_1_120_s_0_350 = 1.70e-11
+ mcm2m1f_ca_w_1_120_s_0_420 = 1.01e-04  mcm2m1f_cc_w_1_120_s_0_420 = 5.32e-11  mcm2m1f_cf_w_1_120_s_0_420 = 1.97e-11
+ mcm2m1f_ca_w_1_120_s_0_560 = 1.01e-04  mcm2m1f_cc_w_1_120_s_0_560 = 4.02e-11  mcm2m1f_cf_w_1_120_s_0_560 = 2.46e-11
+ mcm2m1f_ca_w_1_120_s_0_840 = 1.01e-04  mcm2m1f_cc_w_1_120_s_0_840 = 2.49e-11  mcm2m1f_cf_w_1_120_s_0_840 = 3.26e-11
+ mcm2m1f_ca_w_1_120_s_1_540 = 1.01e-04  mcm2m1f_cc_w_1_120_s_1_540 = 9.15e-12  mcm2m1f_cf_w_1_120_s_1_540 = 4.42e-11
+ mcm2m1f_ca_w_1_120_s_3_500 = 1.01e-04  mcm2m1f_cc_w_1_120_s_3_500 = 8.00e-13  mcm2m1f_cf_w_1_120_s_3_500 = 5.21e-11
+ mcm2m1d_ca_w_0_140_s_0_140 = 1.07e-04  mcm2m1d_cc_w_0_140_s_0_140 = 7.90e-11  mcm2m1d_cf_w_0_140_s_0_140 = 8.48e-12
+ mcm2m1d_ca_w_0_140_s_0_175 = 1.07e-04  mcm2m1d_cc_w_0_140_s_0_175 = 7.71e-11  mcm2m1d_cf_w_0_140_s_0_175 = 1.01e-11
+ mcm2m1d_ca_w_0_140_s_0_210 = 1.07e-04  mcm2m1d_cc_w_0_140_s_0_210 = 7.32e-11  mcm2m1d_cf_w_0_140_s_0_210 = 1.18e-11
+ mcm2m1d_ca_w_0_140_s_0_280 = 1.07e-04  mcm2m1d_cc_w_0_140_s_0_280 = 6.37e-11  mcm2m1d_cf_w_0_140_s_0_280 = 1.49e-11
+ mcm2m1d_ca_w_0_140_s_0_350 = 1.07e-04  mcm2m1d_cc_w_0_140_s_0_350 = 5.39e-11  mcm2m1d_cf_w_0_140_s_0_350 = 1.80e-11
+ mcm2m1d_ca_w_0_140_s_0_420 = 1.07e-04  mcm2m1d_cc_w_0_140_s_0_420 = 4.55e-11  mcm2m1d_cf_w_0_140_s_0_420 = 2.09e-11
+ mcm2m1d_ca_w_0_140_s_0_560 = 1.07e-04  mcm2m1d_cc_w_0_140_s_0_560 = 3.36e-11  mcm2m1d_cf_w_0_140_s_0_560 = 2.60e-11
+ mcm2m1d_ca_w_0_140_s_0_840 = 1.07e-04  mcm2m1d_cc_w_0_140_s_0_840 = 1.98e-11  mcm2m1d_cf_w_0_140_s_0_840 = 3.40e-11
+ mcm2m1d_ca_w_0_140_s_1_540 = 1.07e-04  mcm2m1d_cc_w_0_140_s_1_540 = 6.25e-12  mcm2m1d_cf_w_0_140_s_1_540 = 4.49e-11
+ mcm2m1d_ca_w_0_140_s_3_500 = 1.07e-04  mcm2m1d_cc_w_0_140_s_3_500 = 3.85e-13  mcm2m1d_cf_w_0_140_s_3_500 = 5.06e-11
+ mcm2m1d_ca_w_1_120_s_0_140 = 1.07e-04  mcm2m1d_cc_w_1_120_s_0_140 = 8.95e-11  mcm2m1d_cf_w_1_120_s_0_140 = 8.54e-12
+ mcm2m1d_ca_w_1_120_s_0_175 = 1.07e-04  mcm2m1d_cc_w_1_120_s_0_175 = 8.66e-11  mcm2m1d_cf_w_1_120_s_0_175 = 1.02e-11
+ mcm2m1d_ca_w_1_120_s_0_210 = 1.07e-04  mcm2m1d_cc_w_1_120_s_0_210 = 8.15e-11  mcm2m1d_cf_w_1_120_s_0_210 = 1.19e-11
+ mcm2m1d_ca_w_1_120_s_0_280 = 1.07e-04  mcm2m1d_cc_w_1_120_s_0_280 = 7.06e-11  mcm2m1d_cf_w_1_120_s_0_280 = 1.51e-11
+ mcm2m1d_ca_w_1_120_s_0_350 = 1.07e-04  mcm2m1d_cc_w_1_120_s_0_350 = 5.98e-11  mcm2m1d_cf_w_1_120_s_0_350 = 1.81e-11
+ mcm2m1d_ca_w_1_120_s_0_420 = 1.07e-04  mcm2m1d_cc_w_1_120_s_0_420 = 5.06e-11  mcm2m1d_cf_w_1_120_s_0_420 = 2.11e-11
+ mcm2m1d_ca_w_1_120_s_0_560 = 1.07e-04  mcm2m1d_cc_w_1_120_s_0_560 = 3.73e-11  mcm2m1d_cf_w_1_120_s_0_560 = 2.63e-11
+ mcm2m1d_ca_w_1_120_s_0_840 = 1.07e-04  mcm2m1d_cc_w_1_120_s_0_840 = 2.23e-11  mcm2m1d_cf_w_1_120_s_0_840 = 3.46e-11
+ mcm2m1d_ca_w_1_120_s_1_540 = 1.07e-04  mcm2m1d_cc_w_1_120_s_1_540 = 7.18e-12  mcm2m1d_cf_w_1_120_s_1_540 = 4.62e-11
+ mcm2m1d_ca_w_1_120_s_3_500 = 1.07e-04  mcm2m1d_cc_w_1_120_s_3_500 = 4.20e-13  mcm2m1d_cf_w_1_120_s_3_500 = 5.28e-11
+ mcm2m1p1_ca_w_0_140_s_0_140 = 1.13e-04  mcm2m1p1_cc_w_0_140_s_0_140 = 7.84e-11  mcm2m1p1_cf_w_0_140_s_0_140 = 8.95e-12
+ mcm2m1p1_ca_w_0_140_s_0_175 = 1.13e-04  mcm2m1p1_cc_w_0_140_s_0_175 = 7.64e-11  mcm2m1p1_cf_w_0_140_s_0_175 = 1.07e-11
+ mcm2m1p1_ca_w_0_140_s_0_210 = 1.13e-04  mcm2m1p1_cc_w_0_140_s_0_210 = 7.24e-11  mcm2m1p1_cf_w_0_140_s_0_210 = 1.25e-11
+ mcm2m1p1_ca_w_0_140_s_0_280 = 1.13e-04  mcm2m1p1_cc_w_0_140_s_0_280 = 6.27e-11  mcm2m1p1_cf_w_0_140_s_0_280 = 1.58e-11
+ mcm2m1p1_ca_w_0_140_s_0_350 = 1.13e-04  mcm2m1p1_cc_w_0_140_s_0_350 = 5.28e-11  mcm2m1p1_cf_w_0_140_s_0_350 = 1.91e-11
+ mcm2m1p1_ca_w_0_140_s_0_420 = 1.13e-04  mcm2m1p1_cc_w_0_140_s_0_420 = 4.44e-11  mcm2m1p1_cf_w_0_140_s_0_420 = 2.21e-11
+ mcm2m1p1_ca_w_0_140_s_0_560 = 1.13e-04  mcm2m1p1_cc_w_0_140_s_0_560 = 3.23e-11  mcm2m1p1_cf_w_0_140_s_0_560 = 2.74e-11
+ mcm2m1p1_ca_w_0_140_s_0_840 = 1.13e-04  mcm2m1p1_cc_w_0_140_s_0_840 = 1.84e-11  mcm2m1p1_cf_w_0_140_s_0_840 = 3.58e-11
+ mcm2m1p1_ca_w_0_140_s_1_540 = 1.13e-04  mcm2m1p1_cc_w_0_140_s_1_540 = 5.27e-12  mcm2m1p1_cf_w_0_140_s_1_540 = 4.66e-11
+ mcm2m1p1_ca_w_0_140_s_3_500 = 1.13e-04  mcm2m1p1_cc_w_0_140_s_3_500 = 2.50e-13  mcm2m1p1_cf_w_0_140_s_3_500 = 5.17e-11
+ mcm2m1p1_ca_w_1_120_s_0_140 = 1.13e-04  mcm2m1p1_cc_w_1_120_s_0_140 = 8.76e-11  mcm2m1p1_cf_w_1_120_s_0_140 = 9.06e-12
+ mcm2m1p1_ca_w_1_120_s_0_175 = 1.13e-04  mcm2m1p1_cc_w_1_120_s_0_175 = 8.47e-11  mcm2m1p1_cf_w_1_120_s_0_175 = 1.08e-11
+ mcm2m1p1_ca_w_1_120_s_0_210 = 1.13e-04  mcm2m1p1_cc_w_1_120_s_0_210 = 7.97e-11  mcm2m1p1_cf_w_1_120_s_0_210 = 1.25e-11
+ mcm2m1p1_ca_w_1_120_s_0_280 = 1.13e-04  mcm2m1p1_cc_w_1_120_s_0_280 = 6.85e-11  mcm2m1p1_cf_w_1_120_s_0_280 = 1.60e-11
+ mcm2m1p1_ca_w_1_120_s_0_350 = 1.13e-04  mcm2m1p1_cc_w_1_120_s_0_350 = 5.77e-11  mcm2m1p1_cf_w_1_120_s_0_350 = 1.92e-11
+ mcm2m1p1_ca_w_1_120_s_0_420 = 1.13e-04  mcm2m1p1_cc_w_1_120_s_0_420 = 4.84e-11  mcm2m1p1_cf_w_1_120_s_0_420 = 2.23e-11
+ mcm2m1p1_ca_w_1_120_s_0_560 = 1.13e-04  mcm2m1p1_cc_w_1_120_s_0_560 = 3.54e-11  mcm2m1p1_cf_w_1_120_s_0_560 = 2.77e-11
+ mcm2m1p1_ca_w_1_120_s_0_840 = 1.13e-04  mcm2m1p1_cc_w_1_120_s_0_840 = 2.03e-11  mcm2m1p1_cf_w_1_120_s_0_840 = 3.64e-11
+ mcm2m1p1_ca_w_1_120_s_1_540 = 1.13e-04  mcm2m1p1_cc_w_1_120_s_1_540 = 5.92e-12  mcm2m1p1_cf_w_1_120_s_1_540 = 4.78e-11
+ mcm2m1p1_ca_w_1_120_s_3_500 = 1.13e-04  mcm2m1p1_cc_w_1_120_s_3_500 = 2.95e-13  mcm2m1p1_cf_w_1_120_s_3_500 = 5.36e-11
+ mcm2m1l1_ca_w_0_140_s_0_140 = 1.58e-04  mcm2m1l1_cc_w_0_140_s_0_140 = 7.34e-11  mcm2m1l1_cf_w_0_140_s_0_140 = 1.24e-11
+ mcm2m1l1_ca_w_0_140_s_0_175 = 1.58e-04  mcm2m1l1_cc_w_0_140_s_0_175 = 7.16e-11  mcm2m1l1_cf_w_0_140_s_0_175 = 1.50e-11
+ mcm2m1l1_ca_w_0_140_s_0_210 = 1.58e-04  mcm2m1l1_cc_w_0_140_s_0_210 = 6.69e-11  mcm2m1l1_cf_w_0_140_s_0_210 = 1.75e-11
+ mcm2m1l1_ca_w_0_140_s_0_280 = 1.58e-04  mcm2m1l1_cc_w_0_140_s_0_280 = 5.66e-11  mcm2m1l1_cf_w_0_140_s_0_280 = 2.22e-11
+ mcm2m1l1_ca_w_0_140_s_0_350 = 1.58e-04  mcm2m1l1_cc_w_0_140_s_0_350 = 4.62e-11  mcm2m1l1_cf_w_0_140_s_0_350 = 2.66e-11
+ mcm2m1l1_ca_w_0_140_s_0_420 = 1.58e-04  mcm2m1l1_cc_w_0_140_s_0_420 = 3.76e-11  mcm2m1l1_cf_w_0_140_s_0_420 = 3.07e-11
+ mcm2m1l1_ca_w_0_140_s_0_560 = 1.58e-04  mcm2m1l1_cc_w_0_140_s_0_560 = 2.53e-11  mcm2m1l1_cf_w_0_140_s_0_560 = 3.76e-11
+ mcm2m1l1_ca_w_0_140_s_0_840 = 1.58e-04  mcm2m1l1_cc_w_0_140_s_0_840 = 1.20e-11  mcm2m1l1_cf_w_0_140_s_0_840 = 4.75e-11
+ mcm2m1l1_ca_w_0_140_s_1_540 = 1.58e-04  mcm2m1l1_cc_w_0_140_s_1_540 = 2.00e-12  mcm2m1l1_cf_w_0_140_s_1_540 = 5.69e-11
+ mcm2m1l1_ca_w_0_140_s_3_500 = 1.58e-04  mcm2m1l1_cc_w_0_140_s_3_500 = 3.50e-14  mcm2m1l1_cf_w_0_140_s_3_500 = 5.93e-11
+ mcm2m1l1_ca_w_1_120_s_0_140 = 1.58e-04  mcm2m1l1_cc_w_1_120_s_0_140 = 7.80e-11  mcm2m1l1_cf_w_1_120_s_0_140 = 1.25e-11
+ mcm2m1l1_ca_w_1_120_s_0_175 = 1.58e-04  mcm2m1l1_cc_w_1_120_s_0_175 = 7.49e-11  mcm2m1l1_cf_w_1_120_s_0_175 = 1.51e-11
+ mcm2m1l1_ca_w_1_120_s_0_210 = 1.58e-04  mcm2m1l1_cc_w_1_120_s_0_210 = 7.02e-11  mcm2m1l1_cf_w_1_120_s_0_210 = 1.75e-11
+ mcm2m1l1_ca_w_1_120_s_0_280 = 1.58e-04  mcm2m1l1_cc_w_1_120_s_0_280 = 5.88e-11  mcm2m1l1_cf_w_1_120_s_0_280 = 2.23e-11
+ mcm2m1l1_ca_w_1_120_s_0_350 = 1.58e-04  mcm2m1l1_cc_w_1_120_s_0_350 = 4.80e-11  mcm2m1l1_cf_w_1_120_s_0_350 = 2.68e-11
+ mcm2m1l1_ca_w_1_120_s_0_420 = 1.58e-04  mcm2m1l1_cc_w_1_120_s_0_420 = 3.92e-11  mcm2m1l1_cf_w_1_120_s_0_420 = 3.09e-11
+ mcm2m1l1_ca_w_1_120_s_0_560 = 1.58e-04  mcm2m1l1_cc_w_1_120_s_0_560 = 2.62e-11  mcm2m1l1_cf_w_1_120_s_0_560 = 3.80e-11
+ mcm2m1l1_ca_w_1_120_s_0_840 = 1.58e-04  mcm2m1l1_cc_w_1_120_s_0_840 = 1.24e-11  mcm2m1l1_cf_w_1_120_s_0_840 = 4.81e-11
+ mcm2m1l1_ca_w_1_120_s_1_540 = 1.58e-04  mcm2m1l1_cc_w_1_120_s_1_540 = 2.10e-12  mcm2m1l1_cf_w_1_120_s_1_540 = 5.78e-11
+ mcm2m1l1_ca_w_1_120_s_3_500 = 1.58e-04  mcm2m1l1_cc_w_1_120_s_3_500 = 5.00e-14  mcm2m1l1_cf_w_1_120_s_3_500 = 6.02e-11
+ mcm3m1f_ca_w_0_140_s_0_140 = 4.60e-05  mcm3m1f_cc_w_0_140_s_0_140 = 8.49e-11  mcm3m1f_cf_w_0_140_s_0_140 = 3.84e-12
+ mcm3m1f_ca_w_0_140_s_0_175 = 4.60e-05  mcm3m1f_cc_w_0_140_s_0_175 = 8.40e-11  mcm3m1f_cf_w_0_140_s_0_175 = 4.62e-12
+ mcm3m1f_ca_w_0_140_s_0_210 = 4.60e-05  mcm3m1f_cc_w_0_140_s_0_210 = 8.04e-11  mcm3m1f_cf_w_0_140_s_0_210 = 5.44e-12
+ mcm3m1f_ca_w_0_140_s_0_280 = 4.60e-05  mcm3m1f_cc_w_0_140_s_0_280 = 7.19e-11  mcm3m1f_cf_w_0_140_s_0_280 = 6.93e-12
+ mcm3m1f_ca_w_0_140_s_0_350 = 4.60e-05  mcm3m1f_cc_w_0_140_s_0_350 = 6.26e-11  mcm3m1f_cf_w_0_140_s_0_350 = 8.40e-12
+ mcm3m1f_ca_w_0_140_s_0_420 = 4.60e-05  mcm3m1f_cc_w_0_140_s_0_420 = 5.50e-11  mcm3m1f_cf_w_0_140_s_0_420 = 9.94e-12
+ mcm3m1f_ca_w_0_140_s_0_560 = 4.60e-05  mcm3m1f_cc_w_0_140_s_0_560 = 4.38e-11  mcm3m1f_cf_w_0_140_s_0_560 = 1.27e-11
+ mcm3m1f_ca_w_0_140_s_0_840 = 4.60e-05  mcm3m1f_cc_w_0_140_s_0_840 = 3.02e-11  mcm3m1f_cf_w_0_140_s_0_840 = 1.77e-11
+ mcm3m1f_ca_w_0_140_s_1_540 = 4.60e-05  mcm3m1f_cc_w_0_140_s_1_540 = 1.41e-11  mcm3m1f_cf_w_0_140_s_1_540 = 2.69e-11
+ mcm3m1f_ca_w_0_140_s_3_500 = 4.60e-05  mcm3m1f_cc_w_0_140_s_3_500 = 2.26e-12  mcm3m1f_cf_w_0_140_s_3_500 = 3.68e-11
+ mcm3m1f_ca_w_1_120_s_0_140 = 4.60e-05  mcm3m1f_cc_w_1_120_s_0_140 = 1.04e-10  mcm3m1f_cf_w_1_120_s_0_140 = 3.88e-12
+ mcm3m1f_ca_w_1_120_s_0_175 = 4.60e-05  mcm3m1f_cc_w_1_120_s_0_175 = 1.01e-10  mcm3m1f_cf_w_1_120_s_0_175 = 4.66e-12
+ mcm3m1f_ca_w_1_120_s_0_210 = 4.60e-05  mcm3m1f_cc_w_1_120_s_0_210 = 9.60e-11  mcm3m1f_cf_w_1_120_s_0_210 = 5.44e-12
+ mcm3m1f_ca_w_1_120_s_0_280 = 4.60e-05  mcm3m1f_cc_w_1_120_s_0_280 = 8.52e-11  mcm3m1f_cf_w_1_120_s_0_280 = 6.98e-12
+ mcm3m1f_ca_w_1_120_s_0_350 = 4.60e-05  mcm3m1f_cc_w_1_120_s_0_350 = 7.40e-11  mcm3m1f_cf_w_1_120_s_0_350 = 8.49e-12
+ mcm3m1f_ca_w_1_120_s_0_420 = 4.60e-05  mcm3m1f_cc_w_1_120_s_0_420 = 6.51e-11  mcm3m1f_cf_w_1_120_s_0_420 = 9.97e-12
+ mcm3m1f_ca_w_1_120_s_0_560 = 4.60e-05  mcm3m1f_cc_w_1_120_s_0_560 = 5.18e-11  mcm3m1f_cf_w_1_120_s_0_560 = 1.28e-11
+ mcm3m1f_ca_w_1_120_s_0_840 = 4.60e-05  mcm3m1f_cc_w_1_120_s_0_840 = 3.57e-11  mcm3m1f_cf_w_1_120_s_0_840 = 1.80e-11
+ mcm3m1f_ca_w_1_120_s_1_540 = 4.60e-05  mcm3m1f_cc_w_1_120_s_1_540 = 1.69e-11  mcm3m1f_cf_w_1_120_s_1_540 = 2.79e-11
+ mcm3m1f_ca_w_1_120_s_3_500 = 4.60e-05  mcm3m1f_cc_w_1_120_s_3_500 = 2.78e-12  mcm3m1f_cf_w_1_120_s_3_500 = 3.94e-11
+ mcm3m1d_ca_w_0_140_s_0_140 = 5.25e-05  mcm3m1d_cc_w_0_140_s_0_140 = 8.38e-11  mcm3m1d_cf_w_0_140_s_0_140 = 4.38e-12
+ mcm3m1d_ca_w_0_140_s_0_175 = 5.25e-05  mcm3m1d_cc_w_0_140_s_0_175 = 8.32e-11  mcm3m1d_cf_w_0_140_s_0_175 = 5.27e-12
+ mcm3m1d_ca_w_0_140_s_0_210 = 5.25e-05  mcm3m1d_cc_w_0_140_s_0_210 = 7.96e-11  mcm3m1d_cf_w_0_140_s_0_210 = 6.20e-12
+ mcm3m1d_ca_w_0_140_s_0_280 = 5.25e-05  mcm3m1d_cc_w_0_140_s_0_280 = 7.07e-11  mcm3m1d_cf_w_0_140_s_0_280 = 7.91e-12
+ mcm3m1d_ca_w_0_140_s_0_350 = 5.25e-05  mcm3m1d_cc_w_0_140_s_0_350 = 6.14e-11  mcm3m1d_cf_w_0_140_s_0_350 = 9.59e-12
+ mcm3m1d_ca_w_0_140_s_0_420 = 5.25e-05  mcm3m1d_cc_w_0_140_s_0_420 = 5.36e-11  mcm3m1d_cf_w_0_140_s_0_420 = 1.13e-11
+ mcm3m1d_ca_w_0_140_s_0_560 = 5.25e-05  mcm3m1d_cc_w_0_140_s_0_560 = 4.22e-11  mcm3m1d_cf_w_0_140_s_0_560 = 1.45e-11
+ mcm3m1d_ca_w_0_140_s_0_840 = 5.25e-05  mcm3m1d_cc_w_0_140_s_0_840 = 2.83e-11  mcm3m1d_cf_w_0_140_s_0_840 = 2.00e-11
+ mcm3m1d_ca_w_0_140_s_1_540 = 5.25e-05  mcm3m1d_cc_w_0_140_s_1_540 = 1.24e-11  mcm3m1d_cf_w_0_140_s_1_540 = 2.98e-11
+ mcm3m1d_ca_w_0_140_s_3_500 = 5.25e-05  mcm3m1d_cc_w_0_140_s_3_500 = 1.57e-12  mcm3m1d_cf_w_0_140_s_3_500 = 3.92e-11
+ mcm3m1d_ca_w_1_120_s_0_140 = 5.25e-05  mcm3m1d_cc_w_1_120_s_0_140 = 1.01e-10  mcm3m1d_cf_w_1_120_s_0_140 = 4.44e-12
+ mcm3m1d_ca_w_1_120_s_0_175 = 5.25e-05  mcm3m1d_cc_w_1_120_s_0_175 = 9.82e-11  mcm3m1d_cf_w_1_120_s_0_175 = 5.33e-12
+ mcm3m1d_ca_w_1_120_s_0_210 = 5.25e-05  mcm3m1d_cc_w_1_120_s_0_210 = 9.31e-11  mcm3m1d_cf_w_1_120_s_0_210 = 6.20e-12
+ mcm3m1d_ca_w_1_120_s_0_280 = 5.25e-05  mcm3m1d_cc_w_1_120_s_0_280 = 8.25e-11  mcm3m1d_cf_w_1_120_s_0_280 = 7.95e-12
+ mcm3m1d_ca_w_1_120_s_0_350 = 5.25e-05  mcm3m1d_cc_w_1_120_s_0_350 = 7.14e-11  mcm3m1d_cf_w_1_120_s_0_350 = 9.69e-12
+ mcm3m1d_ca_w_1_120_s_0_420 = 5.25e-05  mcm3m1d_cc_w_1_120_s_0_420 = 6.25e-11  mcm3m1d_cf_w_1_120_s_0_420 = 1.13e-11
+ mcm3m1d_ca_w_1_120_s_0_560 = 5.25e-05  mcm3m1d_cc_w_1_120_s_0_560 = 4.90e-11  mcm3m1d_cf_w_1_120_s_0_560 = 1.46e-11
+ mcm3m1d_ca_w_1_120_s_0_840 = 5.25e-05  mcm3m1d_cc_w_1_120_s_0_840 = 3.28e-11  mcm3m1d_cf_w_1_120_s_0_840 = 2.03e-11
+ mcm3m1d_ca_w_1_120_s_1_540 = 5.25e-05  mcm3m1d_cc_w_1_120_s_1_540 = 1.45e-11  mcm3m1d_cf_w_1_120_s_1_540 = 3.09e-11
+ mcm3m1d_ca_w_1_120_s_3_500 = 5.25e-05  mcm3m1d_cc_w_1_120_s_3_500 = 1.89e-12  mcm3m1d_cf_w_1_120_s_3_500 = 4.17e-11
+ mcm3m1p1_ca_w_0_140_s_0_140 = 5.81e-05  mcm3m1p1_cc_w_0_140_s_0_140 = 8.31e-11  mcm3m1p1_cf_w_0_140_s_0_140 = 4.86e-12
+ mcm3m1p1_ca_w_0_140_s_0_175 = 5.81e-05  mcm3m1p1_cc_w_0_140_s_0_175 = 8.21e-11  mcm3m1p1_cf_w_0_140_s_0_175 = 5.84e-12
+ mcm3m1p1_ca_w_0_140_s_0_210 = 5.81e-05  mcm3m1p1_cc_w_0_140_s_0_210 = 7.89e-11  mcm3m1p1_cf_w_0_140_s_0_210 = 6.87e-12
+ mcm3m1p1_ca_w_0_140_s_0_280 = 5.81e-05  mcm3m1p1_cc_w_0_140_s_0_280 = 6.98e-11  mcm3m1p1_cf_w_0_140_s_0_280 = 8.76e-12
+ mcm3m1p1_ca_w_0_140_s_0_350 = 5.81e-05  mcm3m1p1_cc_w_0_140_s_0_350 = 6.04e-11  mcm3m1p1_cf_w_0_140_s_0_350 = 1.06e-11
+ mcm3m1p1_ca_w_0_140_s_0_420 = 5.81e-05  mcm3m1p1_cc_w_0_140_s_0_420 = 5.20e-11  mcm3m1p1_cf_w_0_140_s_0_420 = 1.25e-11
+ mcm3m1p1_ca_w_0_140_s_0_560 = 5.81e-05  mcm3m1p1_cc_w_0_140_s_0_560 = 4.08e-11  mcm3m1p1_cf_w_0_140_s_0_560 = 1.59e-11
+ mcm3m1p1_ca_w_0_140_s_0_840 = 5.81e-05  mcm3m1p1_cc_w_0_140_s_0_840 = 2.68e-11  mcm3m1p1_cf_w_0_140_s_0_840 = 2.19e-11
+ mcm3m1p1_ca_w_0_140_s_1_540 = 5.81e-05  mcm3m1p1_cc_w_0_140_s_1_540 = 1.10e-11  mcm3m1p1_cf_w_0_140_s_1_540 = 3.22e-11
+ mcm3m1p1_ca_w_0_140_s_3_500 = 5.81e-05  mcm3m1p1_cc_w_0_140_s_3_500 = 1.19e-12  mcm3m1p1_cf_w_0_140_s_3_500 = 4.10e-11
+ mcm3m1p1_ca_w_1_120_s_0_140 = 5.81e-05  mcm3m1p1_cc_w_1_120_s_0_140 = 9.92e-11  mcm3m1p1_cf_w_1_120_s_0_140 = 4.94e-12
+ mcm3m1p1_ca_w_1_120_s_0_175 = 5.81e-05  mcm3m1p1_cc_w_1_120_s_0_175 = 9.62e-11  mcm3m1p1_cf_w_1_120_s_0_175 = 5.93e-12
+ mcm3m1p1_ca_w_1_120_s_0_210 = 5.81e-05  mcm3m1p1_cc_w_1_120_s_0_210 = 9.16e-11  mcm3m1p1_cf_w_1_120_s_0_210 = 6.91e-12
+ mcm3m1p1_ca_w_1_120_s_0_280 = 5.81e-05  mcm3m1p1_cc_w_1_120_s_0_280 = 8.04e-11  mcm3m1p1_cf_w_1_120_s_0_280 = 8.85e-12
+ mcm3m1p1_ca_w_1_120_s_0_350 = 5.81e-05  mcm3m1p1_cc_w_1_120_s_0_350 = 6.95e-11  mcm3m1p1_cf_w_1_120_s_0_350 = 1.07e-11
+ mcm3m1p1_ca_w_1_120_s_0_420 = 5.81e-05  mcm3m1p1_cc_w_1_120_s_0_420 = 6.01e-11  mcm3m1p1_cf_w_1_120_s_0_420 = 1.26e-11
+ mcm3m1p1_ca_w_1_120_s_0_560 = 5.81e-05  mcm3m1p1_cc_w_1_120_s_0_560 = 4.68e-11  mcm3m1p1_cf_w_1_120_s_0_560 = 1.61e-11
+ mcm3m1p1_ca_w_1_120_s_0_840 = 5.81e-05  mcm3m1p1_cc_w_1_120_s_0_840 = 3.08e-11  mcm3m1p1_cf_w_1_120_s_0_840 = 2.23e-11
+ mcm3m1p1_ca_w_1_120_s_1_540 = 5.81e-05  mcm3m1p1_cc_w_1_120_s_1_540 = 1.29e-11  mcm3m1p1_cf_w_1_120_s_1_540 = 3.33e-11
+ mcm3m1p1_ca_w_1_120_s_3_500 = 5.81e-05  mcm3m1p1_cc_w_1_120_s_3_500 = 1.39e-12  mcm3m1p1_cf_w_1_120_s_3_500 = 4.33e-11
+ mcm3m1l1_ca_w_0_140_s_0_140 = 1.03e-04  mcm3m1l1_cc_w_0_140_s_0_140 = 7.90e-11  mcm3m1l1_cf_w_0_140_s_0_140 = 8.37e-12
+ mcm3m1l1_ca_w_0_140_s_0_175 = 1.03e-04  mcm3m1l1_cc_w_0_140_s_0_175 = 7.73e-11  mcm3m1l1_cf_w_0_140_s_0_175 = 1.01e-11
+ mcm3m1l1_ca_w_0_140_s_0_210 = 1.03e-04  mcm3m1l1_cc_w_0_140_s_0_210 = 7.33e-11  mcm3m1l1_cf_w_0_140_s_0_210 = 1.19e-11
+ mcm3m1l1_ca_w_0_140_s_0_280 = 1.03e-04  mcm3m1l1_cc_w_0_140_s_0_280 = 6.36e-11  mcm3m1l1_cf_w_0_140_s_0_280 = 1.51e-11
+ mcm3m1l1_ca_w_0_140_s_0_350 = 1.03e-04  mcm3m1l1_cc_w_0_140_s_0_350 = 5.38e-11  mcm3m1l1_cf_w_0_140_s_0_350 = 1.82e-11
+ mcm3m1l1_ca_w_0_140_s_0_420 = 1.03e-04  mcm3m1l1_cc_w_0_140_s_0_420 = 4.54e-11  mcm3m1l1_cf_w_0_140_s_0_420 = 2.12e-11
+ mcm3m1l1_ca_w_0_140_s_0_560 = 1.03e-04  mcm3m1l1_cc_w_0_140_s_0_560 = 3.34e-11  mcm3m1l1_cf_w_0_140_s_0_560 = 2.66e-11
+ mcm3m1l1_ca_w_0_140_s_0_840 = 1.03e-04  mcm3m1l1_cc_w_0_140_s_0_840 = 1.96e-11  mcm3m1l1_cf_w_0_140_s_0_840 = 3.49e-11
+ mcm3m1l1_ca_w_0_140_s_1_540 = 1.03e-04  mcm3m1l1_cc_w_0_140_s_1_540 = 6.04e-12  mcm3m1l1_cf_w_0_140_s_1_540 = 4.58e-11
+ mcm3m1l1_ca_w_0_140_s_3_500 = 1.03e-04  mcm3m1l1_cc_w_0_140_s_3_500 = 3.35e-13  mcm3m1l1_cf_w_0_140_s_3_500 = 5.15e-11
+ mcm3m1l1_ca_w_1_120_s_0_140 = 1.03e-04  mcm3m1l1_cc_w_1_120_s_0_140 = 8.92e-11  mcm3m1l1_cf_w_1_120_s_0_140 = 8.46e-12
+ mcm3m1l1_ca_w_1_120_s_0_175 = 1.03e-04  mcm3m1l1_cc_w_1_120_s_0_175 = 8.67e-11  mcm3m1l1_cf_w_1_120_s_0_175 = 1.02e-11
+ mcm3m1l1_ca_w_1_120_s_0_210 = 1.03e-04  mcm3m1l1_cc_w_1_120_s_0_210 = 8.20e-11  mcm3m1l1_cf_w_1_120_s_0_210 = 1.19e-11
+ mcm3m1l1_ca_w_1_120_s_0_280 = 1.03e-04  mcm3m1l1_cc_w_1_120_s_0_280 = 7.07e-11  mcm3m1l1_cf_w_1_120_s_0_280 = 1.52e-11
+ mcm3m1l1_ca_w_1_120_s_0_350 = 1.03e-04  mcm3m1l1_cc_w_1_120_s_0_350 = 5.96e-11  mcm3m1l1_cf_w_1_120_s_0_350 = 1.84e-11
+ mcm3m1l1_ca_w_1_120_s_0_420 = 1.03e-04  mcm3m1l1_cc_w_1_120_s_0_420 = 5.04e-11  mcm3m1l1_cf_w_1_120_s_0_420 = 2.13e-11
+ mcm3m1l1_ca_w_1_120_s_0_560 = 1.03e-04  mcm3m1l1_cc_w_1_120_s_0_560 = 3.74e-11  mcm3m1l1_cf_w_1_120_s_0_560 = 2.68e-11
+ mcm3m1l1_ca_w_1_120_s_0_840 = 1.03e-04  mcm3m1l1_cc_w_1_120_s_0_840 = 2.22e-11  mcm3m1l1_cf_w_1_120_s_0_840 = 3.54e-11
+ mcm3m1l1_ca_w_1_120_s_1_540 = 1.03e-04  mcm3m1l1_cc_w_1_120_s_1_540 = 7.17e-12  mcm3m1l1_cf_w_1_120_s_1_540 = 4.72e-11
+ mcm3m1l1_ca_w_1_120_s_3_500 = 1.03e-04  mcm3m1l1_cc_w_1_120_s_3_500 = 3.95e-13  mcm3m1l1_cf_w_1_120_s_3_500 = 5.37e-11
+ mcm4m1f_ca_w_0_140_s_0_140 = 3.30e-05  mcm4m1f_cc_w_0_140_s_0_140 = 8.65e-11  mcm4m1f_cf_w_0_140_s_0_140 = 2.78e-12
+ mcm4m1f_ca_w_0_140_s_0_175 = 3.30e-05  mcm4m1f_cc_w_0_140_s_0_175 = 8.53e-11  mcm4m1f_cf_w_0_140_s_0_175 = 3.35e-12
+ mcm4m1f_ca_w_0_140_s_0_210 = 3.30e-05  mcm4m1f_cc_w_0_140_s_0_210 = 8.22e-11  mcm4m1f_cf_w_0_140_s_0_210 = 3.95e-12
+ mcm4m1f_ca_w_0_140_s_0_280 = 3.30e-05  mcm4m1f_cc_w_0_140_s_0_280 = 7.42e-11  mcm4m1f_cf_w_0_140_s_0_280 = 5.05e-12
+ mcm4m1f_ca_w_0_140_s_0_350 = 3.30e-05  mcm4m1f_cc_w_0_140_s_0_350 = 6.52e-11  mcm4m1f_cf_w_0_140_s_0_350 = 6.14e-12
+ mcm4m1f_ca_w_0_140_s_0_420 = 3.30e-05  mcm4m1f_cc_w_0_140_s_0_420 = 5.75e-11  mcm4m1f_cf_w_0_140_s_0_420 = 7.26e-12
+ mcm4m1f_ca_w_0_140_s_0_560 = 3.30e-05  mcm4m1f_cc_w_0_140_s_0_560 = 4.70e-11  mcm4m1f_cf_w_0_140_s_0_560 = 9.36e-12
+ mcm4m1f_ca_w_0_140_s_0_840 = 3.30e-05  mcm4m1f_cc_w_0_140_s_0_840 = 3.41e-11  mcm4m1f_cf_w_0_140_s_0_840 = 1.32e-11
+ mcm4m1f_ca_w_0_140_s_1_540 = 3.30e-05  mcm4m1f_cc_w_0_140_s_1_540 = 1.83e-11  mcm4m1f_cf_w_0_140_s_1_540 = 2.09e-11
+ mcm4m1f_ca_w_0_140_s_3_500 = 3.30e-05  mcm4m1f_cc_w_0_140_s_3_500 = 4.47e-12  mcm4m1f_cf_w_0_140_s_3_500 = 3.14e-11
+ mcm4m1f_ca_w_1_120_s_0_140 = 3.30e-05  mcm4m1f_cc_w_1_120_s_0_140 = 1.09e-10  mcm4m1f_cf_w_1_120_s_0_140 = 2.81e-12
+ mcm4m1f_ca_w_1_120_s_0_175 = 3.30e-05  mcm4m1f_cc_w_1_120_s_0_175 = 1.06e-10  mcm4m1f_cf_w_1_120_s_0_175 = 3.39e-12
+ mcm4m1f_ca_w_1_120_s_0_210 = 3.30e-05  mcm4m1f_cc_w_1_120_s_0_210 = 1.02e-10  mcm4m1f_cf_w_1_120_s_0_210 = 3.95e-12
+ mcm4m1f_ca_w_1_120_s_0_280 = 3.30e-05  mcm4m1f_cc_w_1_120_s_0_280 = 9.09e-11  mcm4m1f_cf_w_1_120_s_0_280 = 5.08e-12
+ mcm4m1f_ca_w_1_120_s_0_350 = 3.30e-05  mcm4m1f_cc_w_1_120_s_0_350 = 8.01e-11  mcm4m1f_cf_w_1_120_s_0_350 = 6.20e-12
+ mcm4m1f_ca_w_1_120_s_0_420 = 3.30e-05  mcm4m1f_cc_w_1_120_s_0_420 = 7.11e-11  mcm4m1f_cf_w_1_120_s_0_420 = 7.28e-12
+ mcm4m1f_ca_w_1_120_s_0_560 = 3.30e-05  mcm4m1f_cc_w_1_120_s_0_560 = 5.78e-11  mcm4m1f_cf_w_1_120_s_0_560 = 9.40e-12
+ mcm4m1f_ca_w_1_120_s_0_840 = 3.30e-05  mcm4m1f_cc_w_1_120_s_0_840 = 4.18e-11  mcm4m1f_cf_w_1_120_s_0_840 = 1.34e-11
+ mcm4m1f_ca_w_1_120_s_1_540 = 3.30e-05  mcm4m1f_cc_w_1_120_s_1_540 = 2.29e-11  mcm4m1f_cf_w_1_120_s_1_540 = 2.16e-11
+ mcm4m1f_ca_w_1_120_s_3_500 = 3.30e-05  mcm4m1f_cc_w_1_120_s_3_500 = 5.78e-12  mcm4m1f_cf_w_1_120_s_3_500 = 3.39e-11
+ mcm4m1d_ca_w_0_140_s_0_140 = 3.94e-05  mcm4m1d_cc_w_0_140_s_0_140 = 8.58e-11  mcm4m1d_cf_w_0_140_s_0_140 = 3.32e-12
+ mcm4m1d_ca_w_0_140_s_0_175 = 3.94e-05  mcm4m1d_cc_w_0_140_s_0_175 = 8.46e-11  mcm4m1d_cf_w_0_140_s_0_175 = 4.00e-12
+ mcm4m1d_ca_w_0_140_s_0_210 = 3.94e-05  mcm4m1d_cc_w_0_140_s_0_210 = 8.13e-11  mcm4m1d_cf_w_0_140_s_0_210 = 4.71e-12
+ mcm4m1d_ca_w_0_140_s_0_280 = 3.94e-05  mcm4m1d_cc_w_0_140_s_0_280 = 7.31e-11  mcm4m1d_cf_w_0_140_s_0_280 = 6.02e-12
+ mcm4m1d_ca_w_0_140_s_0_350 = 3.94e-05  mcm4m1d_cc_w_0_140_s_0_350 = 6.37e-11  mcm4m1d_cf_w_0_140_s_0_350 = 7.31e-12
+ mcm4m1d_ca_w_0_140_s_0_420 = 3.94e-05  mcm4m1d_cc_w_0_140_s_0_420 = 5.62e-11  mcm4m1d_cf_w_0_140_s_0_420 = 8.64e-12
+ mcm4m1d_ca_w_0_140_s_0_560 = 3.94e-05  mcm4m1d_cc_w_0_140_s_0_560 = 4.53e-11  mcm4m1d_cf_w_0_140_s_0_560 = 1.11e-11
+ mcm4m1d_ca_w_0_140_s_0_840 = 3.94e-05  mcm4m1d_cc_w_0_140_s_0_840 = 3.22e-11  mcm4m1d_cf_w_0_140_s_0_840 = 1.55e-11
+ mcm4m1d_ca_w_0_140_s_1_540 = 3.94e-05  mcm4m1d_cc_w_0_140_s_1_540 = 1.63e-11  mcm4m1d_cf_w_0_140_s_1_540 = 2.41e-11
+ mcm4m1d_ca_w_0_140_s_3_500 = 3.94e-05  mcm4m1d_cc_w_0_140_s_3_500 = 3.42e-12  mcm4m1d_cf_w_0_140_s_3_500 = 3.45e-11
+ mcm4m1d_ca_w_1_120_s_0_140 = 3.94e-05  mcm4m1d_cc_w_1_120_s_0_140 = 1.06e-10  mcm4m1d_cf_w_1_120_s_0_140 = 3.38e-12
+ mcm4m1d_ca_w_1_120_s_0_175 = 3.94e-05  mcm4m1d_cc_w_1_120_s_0_175 = 1.04e-10  mcm4m1d_cf_w_1_120_s_0_175 = 4.06e-12
+ mcm4m1d_ca_w_1_120_s_0_210 = 3.94e-05  mcm4m1d_cc_w_1_120_s_0_210 = 9.91e-11  mcm4m1d_cf_w_1_120_s_0_210 = 4.72e-12
+ mcm4m1d_ca_w_1_120_s_0_280 = 3.94e-05  mcm4m1d_cc_w_1_120_s_0_280 = 8.82e-11  mcm4m1d_cf_w_1_120_s_0_280 = 6.06e-12
+ mcm4m1d_ca_w_1_120_s_0_350 = 3.94e-05  mcm4m1d_cc_w_1_120_s_0_350 = 7.74e-11  mcm4m1d_cf_w_1_120_s_0_350 = 7.38e-12
+ mcm4m1d_ca_w_1_120_s_0_420 = 3.94e-05  mcm4m1d_cc_w_1_120_s_0_420 = 6.84e-11  mcm4m1d_cf_w_1_120_s_0_420 = 8.67e-12
+ mcm4m1d_ca_w_1_120_s_0_560 = 3.94e-05  mcm4m1d_cc_w_1_120_s_0_560 = 5.50e-11  mcm4m1d_cf_w_1_120_s_0_560 = 1.12e-11
+ mcm4m1d_ca_w_1_120_s_0_840 = 3.94e-05  mcm4m1d_cc_w_1_120_s_0_840 = 3.90e-11  mcm4m1d_cf_w_1_120_s_0_840 = 1.58e-11
+ mcm4m1d_ca_w_1_120_s_1_540 = 3.94e-05  mcm4m1d_cc_w_1_120_s_1_540 = 2.02e-11  mcm4m1d_cf_w_1_120_s_1_540 = 2.50e-11
+ mcm4m1d_ca_w_1_120_s_3_500 = 3.94e-05  mcm4m1d_cc_w_1_120_s_3_500 = 4.45e-12  mcm4m1d_cf_w_1_120_s_3_500 = 3.71e-11
+ mcm4m1p1_ca_w_0_140_s_0_140 = 4.51e-05  mcm4m1p1_cc_w_0_140_s_0_140 = 8.53e-11  mcm4m1p1_cf_w_0_140_s_0_140 = 3.79e-12
+ mcm4m1p1_ca_w_0_140_s_0_175 = 4.51e-05  mcm4m1p1_cc_w_0_140_s_0_175 = 8.39e-11  mcm4m1p1_cf_w_0_140_s_0_175 = 4.57e-12
+ mcm4m1p1_ca_w_0_140_s_0_210 = 4.51e-05  mcm4m1p1_cc_w_0_140_s_0_210 = 8.06e-11  mcm4m1p1_cf_w_0_140_s_0_210 = 5.38e-12
+ mcm4m1p1_ca_w_0_140_s_0_280 = 4.51e-05  mcm4m1p1_cc_w_0_140_s_0_280 = 7.22e-11  mcm4m1p1_cf_w_0_140_s_0_280 = 6.88e-12
+ mcm4m1p1_ca_w_0_140_s_0_350 = 4.51e-05  mcm4m1p1_cc_w_0_140_s_0_350 = 6.31e-11  mcm4m1p1_cf_w_0_140_s_0_350 = 8.36e-12
+ mcm4m1p1_ca_w_0_140_s_0_420 = 4.51e-05  mcm4m1p1_cc_w_0_140_s_0_420 = 5.49e-11  mcm4m1p1_cf_w_0_140_s_0_420 = 9.84e-12
+ mcm4m1p1_ca_w_0_140_s_0_560 = 4.51e-05  mcm4m1p1_cc_w_0_140_s_0_560 = 4.40e-11  mcm4m1p1_cf_w_0_140_s_0_560 = 1.26e-11
+ mcm4m1p1_ca_w_0_140_s_0_840 = 4.51e-05  mcm4m1p1_cc_w_0_140_s_0_840 = 3.06e-11  mcm4m1p1_cf_w_0_140_s_0_840 = 1.75e-11
+ mcm4m1p1_ca_w_0_140_s_1_540 = 4.51e-05  mcm4m1p1_cc_w_0_140_s_1_540 = 1.49e-11  mcm4m1p1_cf_w_0_140_s_1_540 = 2.67e-11
+ mcm4m1p1_ca_w_0_140_s_3_500 = 4.51e-05  mcm4m1p1_cc_w_0_140_s_3_500 = 2.77e-12  mcm4m1p1_cf_w_0_140_s_3_500 = 3.67e-11
+ mcm4m1p1_ca_w_1_120_s_0_140 = 4.51e-05  mcm4m1p1_cc_w_1_120_s_0_140 = 1.04e-10  mcm4m1p1_cf_w_1_120_s_0_140 = 3.88e-12
+ mcm4m1p1_ca_w_1_120_s_0_175 = 4.51e-05  mcm4m1p1_cc_w_1_120_s_0_175 = 1.02e-10  mcm4m1p1_cf_w_1_120_s_0_175 = 4.67e-12
+ mcm4m1p1_ca_w_1_120_s_0_210 = 4.51e-05  mcm4m1p1_cc_w_1_120_s_0_210 = 9.69e-11  mcm4m1p1_cf_w_1_120_s_0_210 = 5.43e-12
+ mcm4m1p1_ca_w_1_120_s_0_280 = 4.51e-05  mcm4m1p1_cc_w_1_120_s_0_280 = 8.60e-11  mcm4m1p1_cf_w_1_120_s_0_280 = 6.97e-12
+ mcm4m1p1_ca_w_1_120_s_0_350 = 4.51e-05  mcm4m1p1_cc_w_1_120_s_0_350 = 7.52e-11  mcm4m1p1_cf_w_1_120_s_0_350 = 8.46e-12
+ mcm4m1p1_ca_w_1_120_s_0_420 = 4.51e-05  mcm4m1p1_cc_w_1_120_s_0_420 = 6.61e-11  mcm4m1p1_cf_w_1_120_s_0_420 = 9.92e-12
+ mcm4m1p1_ca_w_1_120_s_0_560 = 4.51e-05  mcm4m1p1_cc_w_1_120_s_0_560 = 5.29e-11  mcm4m1p1_cf_w_1_120_s_0_560 = 1.27e-11
+ mcm4m1p1_ca_w_1_120_s_0_840 = 4.51e-05  mcm4m1p1_cc_w_1_120_s_0_840 = 3.69e-11  mcm4m1p1_cf_w_1_120_s_0_840 = 1.78e-11
+ mcm4m1p1_ca_w_1_120_s_1_540 = 4.51e-05  mcm4m1p1_cc_w_1_120_s_1_540 = 1.84e-11  mcm4m1p1_cf_w_1_120_s_1_540 = 2.76e-11
+ mcm4m1p1_ca_w_1_120_s_3_500 = 4.51e-05  mcm4m1p1_cc_w_1_120_s_3_500 = 3.63e-12  mcm4m1p1_cf_w_1_120_s_3_500 = 3.95e-11
+ mcm4m1l1_ca_w_0_140_s_0_140 = 9.00e-05  mcm4m1l1_cc_w_0_140_s_0_140 = 8.06e-11  mcm4m1l1_cf_w_0_140_s_0_140 = 7.31e-12
+ mcm4m1l1_ca_w_0_140_s_0_175 = 9.00e-05  mcm4m1l1_cc_w_0_140_s_0_175 = 7.90e-11  mcm4m1l1_cf_w_0_140_s_0_175 = 8.88e-12
+ mcm4m1l1_ca_w_0_140_s_0_210 = 9.00e-05  mcm4m1l1_cc_w_0_140_s_0_210 = 7.50e-11  mcm4m1l1_cf_w_0_140_s_0_210 = 1.04e-11
+ mcm4m1l1_ca_w_0_140_s_0_280 = 9.00e-05  mcm4m1l1_cc_w_0_140_s_0_280 = 6.60e-11  mcm4m1l1_cf_w_0_140_s_0_280 = 1.33e-11
+ mcm4m1l1_ca_w_0_140_s_0_350 = 9.00e-05  mcm4m1l1_cc_w_0_140_s_0_350 = 5.58e-11  mcm4m1l1_cf_w_0_140_s_0_350 = 1.60e-11
+ mcm4m1l1_ca_w_0_140_s_0_420 = 9.00e-05  mcm4m1l1_cc_w_0_140_s_0_420 = 4.78e-11  mcm4m1l1_cf_w_0_140_s_0_420 = 1.86e-11
+ mcm4m1l1_ca_w_0_140_s_0_560 = 9.00e-05  mcm4m1l1_cc_w_0_140_s_0_560 = 3.65e-11  mcm4m1l1_cf_w_0_140_s_0_560 = 2.34e-11
+ mcm4m1l1_ca_w_0_140_s_0_840 = 9.00e-05  mcm4m1l1_cc_w_0_140_s_0_840 = 2.30e-11  mcm4m1l1_cf_w_0_140_s_0_840 = 3.09e-11
+ mcm4m1l1_ca_w_0_140_s_1_540 = 9.00e-05  mcm4m1l1_cc_w_0_140_s_1_540 = 8.93e-12  mcm4m1l1_cf_w_0_140_s_1_540 = 4.17e-11
+ mcm4m1l1_ca_w_0_140_s_3_500 = 9.00e-05  mcm4m1l1_cc_w_0_140_s_3_500 = 1.13e-12  mcm4m1l1_cf_w_0_140_s_3_500 = 4.92e-11
+ mcm4m1l1_ca_w_1_120_s_0_140 = 9.00e-05  mcm4m1l1_cc_w_1_120_s_0_140 = 9.50e-11  mcm4m1l1_cf_w_1_120_s_0_140 = 7.40e-12
+ mcm4m1l1_ca_w_1_120_s_0_175 = 9.00e-05  mcm4m1l1_cc_w_1_120_s_0_175 = 9.21e-11  mcm4m1l1_cf_w_1_120_s_0_175 = 8.97e-12
+ mcm4m1l1_ca_w_1_120_s_0_210 = 9.00e-05  mcm4m1l1_cc_w_1_120_s_0_210 = 8.74e-11  mcm4m1l1_cf_w_1_120_s_0_210 = 1.05e-11
+ mcm4m1l1_ca_w_1_120_s_0_280 = 9.00e-05  mcm4m1l1_cc_w_1_120_s_0_280 = 7.64e-11  mcm4m1l1_cf_w_1_120_s_0_280 = 1.34e-11
+ mcm4m1l1_ca_w_1_120_s_0_350 = 9.00e-05  mcm4m1l1_cc_w_1_120_s_0_350 = 6.55e-11  mcm4m1l1_cf_w_1_120_s_0_350 = 1.61e-11
+ mcm4m1l1_ca_w_1_120_s_0_420 = 9.00e-05  mcm4m1l1_cc_w_1_120_s_0_420 = 5.64e-11  mcm4m1l1_cf_w_1_120_s_0_420 = 1.88e-11
+ mcm4m1l1_ca_w_1_120_s_0_560 = 9.00e-05  mcm4m1l1_cc_w_1_120_s_0_560 = 4.33e-11  mcm4m1l1_cf_w_1_120_s_0_560 = 2.34e-11
+ mcm4m1l1_ca_w_1_120_s_0_840 = 9.00e-05  mcm4m1l1_cc_w_1_120_s_0_840 = 2.82e-11  mcm4m1l1_cf_w_1_120_s_0_840 = 3.12e-11
+ mcm4m1l1_ca_w_1_120_s_1_540 = 9.00e-05  mcm4m1l1_cc_w_1_120_s_1_540 = 1.18e-11  mcm4m1l1_cf_w_1_120_s_1_540 = 4.30e-11
+ mcm4m1l1_ca_w_1_120_s_3_500 = 9.00e-05  mcm4m1l1_cc_w_1_120_s_3_500 = 1.71e-12  mcm4m1l1_cf_w_1_120_s_3_500 = 5.24e-11
+ mcm5m1f_ca_w_0_140_s_0_140 = 2.85e-05  mcm5m1f_cc_w_0_140_s_0_140 = 8.70e-11  mcm5m1f_cf_w_0_140_s_0_140 = 2.41e-12
+ mcm5m1f_ca_w_0_140_s_0_175 = 2.85e-05  mcm5m1f_cc_w_0_140_s_0_175 = 8.61e-11  mcm5m1f_cf_w_0_140_s_0_175 = 2.90e-12
+ mcm5m1f_ca_w_0_140_s_0_210 = 2.85e-05  mcm5m1f_cc_w_0_140_s_0_210 = 8.29e-11  mcm5m1f_cf_w_0_140_s_0_210 = 3.42e-12
+ mcm5m1f_ca_w_0_140_s_0_280 = 2.85e-05  mcm5m1f_cc_w_0_140_s_0_280 = 7.50e-11  mcm5m1f_cf_w_0_140_s_0_280 = 4.37e-12
+ mcm5m1f_ca_w_0_140_s_0_350 = 2.85e-05  mcm5m1f_cc_w_0_140_s_0_350 = 6.63e-11  mcm5m1f_cf_w_0_140_s_0_350 = 5.33e-12
+ mcm5m1f_ca_w_0_140_s_0_420 = 2.85e-05  mcm5m1f_cc_w_0_140_s_0_420 = 5.84e-11  mcm5m1f_cf_w_0_140_s_0_420 = 6.30e-12
+ mcm5m1f_ca_w_0_140_s_0_560 = 2.85e-05  mcm5m1f_cc_w_0_140_s_0_560 = 4.81e-11  mcm5m1f_cf_w_0_140_s_0_560 = 8.13e-12
+ mcm5m1f_ca_w_0_140_s_0_840 = 2.85e-05  mcm5m1f_cc_w_0_140_s_0_840 = 3.56e-11  mcm5m1f_cf_w_0_140_s_0_840 = 1.15e-11
+ mcm5m1f_ca_w_0_140_s_1_540 = 2.85e-05  mcm5m1f_cc_w_0_140_s_1_540 = 2.03e-11  mcm5m1f_cf_w_0_140_s_1_540 = 1.85e-11
+ mcm5m1f_ca_w_0_140_s_3_500 = 2.85e-05  mcm5m1f_cc_w_0_140_s_3_500 = 6.02e-12  mcm5m1f_cf_w_0_140_s_3_500 = 2.89e-11
+ mcm5m1f_ca_w_1_120_s_0_140 = 2.85e-05  mcm5m1f_cc_w_1_120_s_0_140 = 1.11e-10  mcm5m1f_cf_w_1_120_s_0_140 = 2.44e-12
+ mcm5m1f_ca_w_1_120_s_0_175 = 2.85e-05  mcm5m1f_cc_w_1_120_s_0_175 = 1.09e-10  mcm5m1f_cf_w_1_120_s_0_175 = 2.93e-12
+ mcm5m1f_ca_w_1_120_s_0_210 = 2.85e-05  mcm5m1f_cc_w_1_120_s_0_210 = 1.04e-10  mcm5m1f_cf_w_1_120_s_0_210 = 3.42e-12
+ mcm5m1f_ca_w_1_120_s_0_280 = 2.85e-05  mcm5m1f_cc_w_1_120_s_0_280 = 9.28e-11  mcm5m1f_cf_w_1_120_s_0_280 = 4.42e-12
+ mcm5m1f_ca_w_1_120_s_0_350 = 2.85e-05  mcm5m1f_cc_w_1_120_s_0_350 = 8.23e-11  mcm5m1f_cf_w_1_120_s_0_350 = 5.37e-12
+ mcm5m1f_ca_w_1_120_s_0_420 = 2.85e-05  mcm5m1f_cc_w_1_120_s_0_420 = 7.34e-11  mcm5m1f_cf_w_1_120_s_0_420 = 6.31e-12
+ mcm5m1f_ca_w_1_120_s_0_560 = 2.85e-05  mcm5m1f_cc_w_1_120_s_0_560 = 6.05e-11  mcm5m1f_cf_w_1_120_s_0_560 = 8.16e-12
+ mcm5m1f_ca_w_1_120_s_0_840 = 2.85e-05  mcm5m1f_cc_w_1_120_s_0_840 = 4.48e-11  mcm5m1f_cf_w_1_120_s_0_840 = 1.17e-11
+ mcm5m1f_ca_w_1_120_s_1_540 = 2.85e-05  mcm5m1f_cc_w_1_120_s_1_540 = 2.60e-11  mcm5m1f_cf_w_1_120_s_1_540 = 1.91e-11
+ mcm5m1f_ca_w_1_120_s_3_500 = 2.85e-05  mcm5m1f_cc_w_1_120_s_3_500 = 8.05e-12  mcm5m1f_cf_w_1_120_s_3_500 = 3.12e-11
+ mcm5m1d_ca_w_0_140_s_0_140 = 3.49e-05  mcm5m1d_cc_w_0_140_s_0_140 = 8.63e-11  mcm5m1d_cf_w_0_140_s_0_140 = 2.94e-12
+ mcm5m1d_ca_w_0_140_s_0_175 = 3.49e-05  mcm5m1d_cc_w_0_140_s_0_175 = 8.52e-11  mcm5m1d_cf_w_0_140_s_0_175 = 3.55e-12
+ mcm5m1d_ca_w_0_140_s_0_210 = 3.49e-05  mcm5m1d_cc_w_0_140_s_0_210 = 8.19e-11  mcm5m1d_cf_w_0_140_s_0_210 = 4.17e-12
+ mcm5m1d_ca_w_0_140_s_0_280 = 3.49e-05  mcm5m1d_cc_w_0_140_s_0_280 = 7.39e-11  mcm5m1d_cf_w_0_140_s_0_280 = 5.35e-12
+ mcm5m1d_ca_w_0_140_s_0_350 = 3.49e-05  mcm5m1d_cc_w_0_140_s_0_350 = 6.50e-11  mcm5m1d_cf_w_0_140_s_0_350 = 6.50e-12
+ mcm5m1d_ca_w_0_140_s_0_420 = 3.49e-05  mcm5m1d_cc_w_0_140_s_0_420 = 5.70e-11  mcm5m1d_cf_w_0_140_s_0_420 = 7.68e-12
+ mcm5m1d_ca_w_0_140_s_0_560 = 3.49e-05  mcm5m1d_cc_w_0_140_s_0_560 = 4.65e-11  mcm5m1d_cf_w_0_140_s_0_560 = 9.88e-12
+ mcm5m1d_ca_w_0_140_s_0_840 = 3.49e-05  mcm5m1d_cc_w_0_140_s_0_840 = 3.37e-11  mcm5m1d_cf_w_0_140_s_0_840 = 1.39e-11
+ mcm5m1d_ca_w_0_140_s_1_540 = 3.49e-05  mcm5m1d_cc_w_0_140_s_1_540 = 1.82e-11  mcm5m1d_cf_w_0_140_s_1_540 = 2.18e-11
+ mcm5m1d_ca_w_0_140_s_3_500 = 3.49e-05  mcm5m1d_cc_w_0_140_s_3_500 = 4.73e-12  mcm5m1d_cf_w_0_140_s_3_500 = 3.23e-11
+ mcm5m1d_ca_w_1_120_s_0_140 = 3.49e-05  mcm5m1d_cc_w_1_120_s_0_140 = 1.08e-10  mcm5m1d_cf_w_1_120_s_0_140 = 3.00e-12
+ mcm5m1d_ca_w_1_120_s_0_175 = 3.49e-05  mcm5m1d_cc_w_1_120_s_0_175 = 1.06e-10  mcm5m1d_cf_w_1_120_s_0_175 = 3.61e-12
+ mcm5m1d_ca_w_1_120_s_0_210 = 3.49e-05  mcm5m1d_cc_w_1_120_s_0_210 = 1.01e-10  mcm5m1d_cf_w_1_120_s_0_210 = 4.19e-12
+ mcm5m1d_ca_w_1_120_s_0_280 = 3.49e-05  mcm5m1d_cc_w_1_120_s_0_280 = 9.02e-11  mcm5m1d_cf_w_1_120_s_0_280 = 5.40e-12
+ mcm5m1d_ca_w_1_120_s_0_350 = 3.49e-05  mcm5m1d_cc_w_1_120_s_0_350 = 7.95e-11  mcm5m1d_cf_w_1_120_s_0_350 = 6.56e-12
+ mcm5m1d_ca_w_1_120_s_0_420 = 3.49e-05  mcm5m1d_cc_w_1_120_s_0_420 = 7.08e-11  mcm5m1d_cf_w_1_120_s_0_420 = 7.71e-12
+ mcm5m1d_ca_w_1_120_s_0_560 = 3.49e-05  mcm5m1d_cc_w_1_120_s_0_560 = 5.77e-11  mcm5m1d_cf_w_1_120_s_0_560 = 9.93e-12
+ mcm5m1d_ca_w_1_120_s_0_840 = 3.49e-05  mcm5m1d_cc_w_1_120_s_0_840 = 4.19e-11  mcm5m1d_cf_w_1_120_s_0_840 = 1.41e-11
+ mcm5m1d_ca_w_1_120_s_1_540 = 3.49e-05  mcm5m1d_cc_w_1_120_s_1_540 = 2.33e-11  mcm5m1d_cf_w_1_120_s_1_540 = 2.25e-11
+ mcm5m1d_ca_w_1_120_s_3_500 = 3.49e-05  mcm5m1d_cc_w_1_120_s_3_500 = 6.47e-12  mcm5m1d_cf_w_1_120_s_3_500 = 3.49e-11
+ mcm5m1p1_ca_w_0_140_s_0_140 = 4.06e-05  mcm5m1p1_cc_w_0_140_s_0_140 = 8.57e-11  mcm5m1p1_cf_w_0_140_s_0_140 = 3.42e-12
+ mcm5m1p1_ca_w_0_140_s_0_175 = 4.06e-05  mcm5m1p1_cc_w_0_140_s_0_175 = 8.45e-11  mcm5m1p1_cf_w_0_140_s_0_175 = 4.12e-12
+ mcm5m1p1_ca_w_0_140_s_0_210 = 4.06e-05  mcm5m1p1_cc_w_0_140_s_0_210 = 8.09e-11  mcm5m1p1_cf_w_0_140_s_0_210 = 4.84e-12
+ mcm5m1p1_ca_w_0_140_s_0_280 = 4.06e-05  mcm5m1p1_cc_w_0_140_s_0_280 = 7.30e-11  mcm5m1p1_cf_w_0_140_s_0_280 = 6.20e-12
+ mcm5m1p1_ca_w_0_140_s_0_350 = 4.06e-05  mcm5m1p1_cc_w_0_140_s_0_350 = 6.40e-11  mcm5m1p1_cf_w_0_140_s_0_350 = 7.54e-12
+ mcm5m1p1_ca_w_0_140_s_0_420 = 4.06e-05  mcm5m1p1_cc_w_0_140_s_0_420 = 5.59e-11  mcm5m1p1_cf_w_0_140_s_0_420 = 8.89e-12
+ mcm5m1p1_ca_w_0_140_s_0_560 = 4.06e-05  mcm5m1p1_cc_w_0_140_s_0_560 = 4.51e-11  mcm5m1p1_cf_w_0_140_s_0_560 = 1.14e-11
+ mcm5m1p1_ca_w_0_140_s_0_840 = 4.06e-05  mcm5m1p1_cc_w_0_140_s_0_840 = 3.22e-11  mcm5m1p1_cf_w_0_140_s_0_840 = 1.58e-11
+ mcm5m1p1_ca_w_0_140_s_1_540 = 4.06e-05  mcm5m1p1_cc_w_0_140_s_1_540 = 1.67e-11  mcm5m1p1_cf_w_0_140_s_1_540 = 2.45e-11
+ mcm5m1p1_ca_w_0_140_s_3_500 = 4.06e-05  mcm5m1p1_cc_w_0_140_s_3_500 = 3.95e-12  mcm5m1p1_cf_w_0_140_s_3_500 = 3.49e-11
+ mcm5m1p1_ca_w_1_120_s_0_140 = 4.06e-05  mcm5m1p1_cc_w_1_120_s_0_140 = 1.07e-10  mcm5m1p1_cf_w_1_120_s_0_140 = 3.51e-12
+ mcm5m1p1_ca_w_1_120_s_0_175 = 4.06e-05  mcm5m1p1_cc_w_1_120_s_0_175 = 1.04e-10  mcm5m1p1_cf_w_1_120_s_0_175 = 4.22e-12
+ mcm5m1p1_ca_w_1_120_s_0_210 = 4.06e-05  mcm5m1p1_cc_w_1_120_s_0_210 = 9.94e-11  mcm5m1p1_cf_w_1_120_s_0_210 = 4.91e-12
+ mcm5m1p1_ca_w_1_120_s_0_280 = 4.06e-05  mcm5m1p1_cc_w_1_120_s_0_280 = 8.81e-11  mcm5m1p1_cf_w_1_120_s_0_280 = 6.31e-12
+ mcm5m1p1_ca_w_1_120_s_0_350 = 4.06e-05  mcm5m1p1_cc_w_1_120_s_0_350 = 7.79e-11  mcm5m1p1_cf_w_1_120_s_0_350 = 7.64e-12
+ mcm5m1p1_ca_w_1_120_s_0_420 = 4.06e-05  mcm5m1p1_cc_w_1_120_s_0_420 = 6.87e-11  mcm5m1p1_cf_w_1_120_s_0_420 = 8.96e-12
+ mcm5m1p1_ca_w_1_120_s_0_560 = 4.06e-05  mcm5m1p1_cc_w_1_120_s_0_560 = 5.56e-11  mcm5m1p1_cf_w_1_120_s_0_560 = 1.15e-11
+ mcm5m1p1_ca_w_1_120_s_0_840 = 4.06e-05  mcm5m1p1_cc_w_1_120_s_0_840 = 3.98e-11  mcm5m1p1_cf_w_1_120_s_0_840 = 1.62e-11
+ mcm5m1p1_ca_w_1_120_s_1_540 = 4.06e-05  mcm5m1p1_cc_w_1_120_s_1_540 = 2.14e-11  mcm5m1p1_cf_w_1_120_s_1_540 = 2.53e-11
+ mcm5m1p1_ca_w_1_120_s_3_500 = 4.06e-05  mcm5m1p1_cc_w_1_120_s_3_500 = 5.51e-12  mcm5m1p1_cf_w_1_120_s_3_500 = 3.76e-11
+ mcm5m1l1_ca_w_0_140_s_0_140 = 8.55e-05  mcm5m1l1_cc_w_0_140_s_0_140 = 8.12e-11  mcm5m1l1_cf_w_0_140_s_0_140 = 6.93e-12
+ mcm5m1l1_ca_w_0_140_s_0_175 = 8.55e-05  mcm5m1l1_cc_w_0_140_s_0_175 = 7.93e-11  mcm5m1l1_cf_w_0_140_s_0_175 = 8.43e-12
+ mcm5m1l1_ca_w_0_140_s_0_210 = 8.55e-05  mcm5m1l1_cc_w_0_140_s_0_210 = 7.56e-11  mcm5m1l1_cf_w_0_140_s_0_210 = 9.87e-12
+ mcm5m1l1_ca_w_0_140_s_0_280 = 8.55e-05  mcm5m1l1_cc_w_0_140_s_0_280 = 6.67e-11  mcm5m1l1_cf_w_0_140_s_0_280 = 1.26e-11
+ mcm5m1l1_ca_w_0_140_s_0_350 = 8.55e-05  mcm5m1l1_cc_w_0_140_s_0_350 = 5.68e-11  mcm5m1l1_cf_w_0_140_s_0_350 = 1.52e-11
+ mcm5m1l1_ca_w_0_140_s_0_420 = 8.55e-05  mcm5m1l1_cc_w_0_140_s_0_420 = 4.91e-11  mcm5m1l1_cf_w_0_140_s_0_420 = 1.77e-11
+ mcm5m1l1_ca_w_0_140_s_0_560 = 8.55e-05  mcm5m1l1_cc_w_0_140_s_0_560 = 3.76e-11  mcm5m1l1_cf_w_0_140_s_0_560 = 2.22e-11
+ mcm5m1l1_ca_w_0_140_s_0_840 = 8.55e-05  mcm5m1l1_cc_w_0_140_s_0_840 = 2.45e-11  mcm5m1l1_cf_w_0_140_s_0_840 = 2.94e-11
+ mcm5m1l1_ca_w_0_140_s_1_540 = 8.55e-05  mcm5m1l1_cc_w_0_140_s_1_540 = 1.03e-11  mcm5m1l1_cf_w_0_140_s_1_540 = 4.01e-11
+ mcm5m1l1_ca_w_0_140_s_3_500 = 8.55e-05  mcm5m1l1_cc_w_0_140_s_3_500 = 1.78e-12  mcm5m1l1_cf_w_0_140_s_3_500 = 4.82e-11
+ mcm5m1l1_ca_w_1_120_s_0_140 = 8.55e-05  mcm5m1l1_cc_w_1_120_s_0_140 = 9.75e-11  mcm5m1l1_cf_w_1_120_s_0_140 = 7.03e-12
+ mcm5m1l1_ca_w_1_120_s_0_175 = 8.55e-05  mcm5m1l1_cc_w_1_120_s_0_175 = 9.44e-11  mcm5m1l1_cf_w_1_120_s_0_175 = 8.51e-12
+ mcm5m1l1_ca_w_1_120_s_0_210 = 8.55e-05  mcm5m1l1_cc_w_1_120_s_0_210 = 8.97e-11  mcm5m1l1_cf_w_1_120_s_0_210 = 9.93e-12
+ mcm5m1l1_ca_w_1_120_s_0_280 = 8.55e-05  mcm5m1l1_cc_w_1_120_s_0_280 = 7.87e-11  mcm5m1l1_cf_w_1_120_s_0_280 = 1.27e-11
+ mcm5m1l1_ca_w_1_120_s_0_350 = 8.55e-05  mcm5m1l1_cc_w_1_120_s_0_350 = 6.78e-11  mcm5m1l1_cf_w_1_120_s_0_350 = 1.53e-11
+ mcm5m1l1_ca_w_1_120_s_0_420 = 8.55e-05  mcm5m1l1_cc_w_1_120_s_0_420 = 5.88e-11  mcm5m1l1_cf_w_1_120_s_0_420 = 1.78e-11
+ mcm5m1l1_ca_w_1_120_s_0_560 = 8.55e-05  mcm5m1l1_cc_w_1_120_s_0_560 = 4.60e-11  mcm5m1l1_cf_w_1_120_s_0_560 = 2.23e-11
+ mcm5m1l1_ca_w_1_120_s_0_840 = 8.55e-05  mcm5m1l1_cc_w_1_120_s_0_840 = 3.09e-11  mcm5m1l1_cf_w_1_120_s_0_840 = 2.97e-11
+ mcm5m1l1_ca_w_1_120_s_1_540 = 8.55e-05  mcm5m1l1_cc_w_1_120_s_1_540 = 1.44e-11  mcm5m1l1_cf_w_1_120_s_1_540 = 4.14e-11
+ mcm5m1l1_ca_w_1_120_s_3_500 = 8.55e-05  mcm5m1l1_cc_w_1_120_s_3_500 = 2.91e-12  mcm5m1l1_cf_w_1_120_s_3_500 = 5.17e-11
+ mcrdlm1f_ca_w_0_140_s_0_140 = 2.27e-05  mcrdlm1f_cc_w_0_140_s_0_140 = 8.78e-11  mcrdlm1f_cf_w_0_140_s_0_140 = 1.92e-12
+ mcrdlm1f_ca_w_0_140_s_0_175 = 2.27e-05  mcrdlm1f_cc_w_0_140_s_0_175 = 8.66e-11  mcrdlm1f_cf_w_0_140_s_0_175 = 2.31e-12
+ mcrdlm1f_ca_w_0_140_s_0_210 = 2.27e-05  mcrdlm1f_cc_w_0_140_s_0_210 = 8.34e-11  mcrdlm1f_cf_w_0_140_s_0_210 = 2.71e-12
+ mcrdlm1f_ca_w_0_140_s_0_280 = 2.27e-05  mcrdlm1f_cc_w_0_140_s_0_280 = 7.61e-11  mcrdlm1f_cf_w_0_140_s_0_280 = 3.48e-12
+ mcrdlm1f_ca_w_0_140_s_0_350 = 2.27e-05  mcrdlm1f_cc_w_0_140_s_0_350 = 6.70e-11  mcrdlm1f_cf_w_0_140_s_0_350 = 4.24e-12
+ mcrdlm1f_ca_w_0_140_s_0_420 = 2.27e-05  mcrdlm1f_cc_w_0_140_s_0_420 = 5.97e-11  mcrdlm1f_cf_w_0_140_s_0_420 = 5.03e-12
+ mcrdlm1f_ca_w_0_140_s_0_560 = 2.27e-05  mcrdlm1f_cc_w_0_140_s_0_560 = 4.97e-11  mcrdlm1f_cf_w_0_140_s_0_560 = 6.47e-12
+ mcrdlm1f_ca_w_0_140_s_0_840 = 2.27e-05  mcrdlm1f_cc_w_0_140_s_0_840 = 3.77e-11  mcrdlm1f_cf_w_0_140_s_0_840 = 9.22e-12
+ mcrdlm1f_ca_w_0_140_s_1_540 = 2.27e-05  mcrdlm1f_cc_w_0_140_s_1_540 = 2.34e-11  mcrdlm1f_cf_w_0_140_s_1_540 = 1.51e-11
+ mcrdlm1f_ca_w_0_140_s_3_500 = 2.27e-05  mcrdlm1f_cc_w_0_140_s_3_500 = 9.18e-12  mcrdlm1f_cf_w_0_140_s_3_500 = 2.49e-11
+ mcrdlm1f_ca_w_1_120_s_0_140 = 2.27e-05  mcrdlm1f_cc_w_1_120_s_0_140 = 1.14e-10  mcrdlm1f_cf_w_1_120_s_0_140 = 1.95e-12
+ mcrdlm1f_ca_w_1_120_s_0_175 = 2.27e-05  mcrdlm1f_cc_w_1_120_s_0_175 = 1.12e-10  mcrdlm1f_cf_w_1_120_s_0_175 = 2.35e-12
+ mcrdlm1f_ca_w_1_120_s_0_210 = 2.27e-05  mcrdlm1f_cc_w_1_120_s_0_210 = 1.07e-10  mcrdlm1f_cf_w_1_120_s_0_210 = 2.73e-12
+ mcrdlm1f_ca_w_1_120_s_0_280 = 2.27e-05  mcrdlm1f_cc_w_1_120_s_0_280 = 9.58e-11  mcrdlm1f_cf_w_1_120_s_0_280 = 3.52e-12
+ mcrdlm1f_ca_w_1_120_s_0_350 = 2.27e-05  mcrdlm1f_cc_w_1_120_s_0_350 = 8.59e-11  mcrdlm1f_cf_w_1_120_s_0_350 = 4.29e-12
+ mcrdlm1f_ca_w_1_120_s_0_420 = 2.27e-05  mcrdlm1f_cc_w_1_120_s_0_420 = 7.69e-11  mcrdlm1f_cf_w_1_120_s_0_420 = 5.05e-12
+ mcrdlm1f_ca_w_1_120_s_0_560 = 2.27e-05  mcrdlm1f_cc_w_1_120_s_0_560 = 6.44e-11  mcrdlm1f_cf_w_1_120_s_0_560 = 6.51e-12
+ mcrdlm1f_ca_w_1_120_s_0_840 = 2.27e-05  mcrdlm1f_cc_w_1_120_s_0_840 = 4.92e-11  mcrdlm1f_cf_w_1_120_s_0_840 = 9.33e-12
+ mcrdlm1f_ca_w_1_120_s_1_540 = 2.27e-05  mcrdlm1f_cc_w_1_120_s_1_540 = 3.12e-11  mcrdlm1f_cf_w_1_120_s_1_540 = 1.55e-11
+ mcrdlm1f_ca_w_1_120_s_3_500 = 2.27e-05  mcrdlm1f_cc_w_1_120_s_3_500 = 1.31e-11  mcrdlm1f_cf_w_1_120_s_3_500 = 2.68e-11
+ mcrdlm1d_ca_w_0_140_s_0_140 = 2.91e-05  mcrdlm1d_cc_w_0_140_s_0_140 = 8.71e-11  mcrdlm1d_cf_w_0_140_s_0_140 = 2.45e-12
+ mcrdlm1d_ca_w_0_140_s_0_175 = 2.91e-05  mcrdlm1d_cc_w_0_140_s_0_175 = 8.55e-11  mcrdlm1d_cf_w_0_140_s_0_175 = 2.96e-12
+ mcrdlm1d_ca_w_0_140_s_0_210 = 2.91e-05  mcrdlm1d_cc_w_0_140_s_0_210 = 8.25e-11  mcrdlm1d_cf_w_0_140_s_0_210 = 3.47e-12
+ mcrdlm1d_ca_w_0_140_s_0_280 = 2.91e-05  mcrdlm1d_cc_w_0_140_s_0_280 = 7.48e-11  mcrdlm1d_cf_w_0_140_s_0_280 = 4.46e-12
+ mcrdlm1d_ca_w_0_140_s_0_350 = 2.91e-05  mcrdlm1d_cc_w_0_140_s_0_350 = 6.58e-11  mcrdlm1d_cf_w_0_140_s_0_350 = 5.42e-12
+ mcrdlm1d_ca_w_0_140_s_0_420 = 2.91e-05  mcrdlm1d_cc_w_0_140_s_0_420 = 5.84e-11  mcrdlm1d_cf_w_0_140_s_0_420 = 6.41e-12
+ mcrdlm1d_ca_w_0_140_s_0_560 = 2.91e-05  mcrdlm1d_cc_w_0_140_s_0_560 = 4.81e-11  mcrdlm1d_cf_w_0_140_s_0_560 = 8.23e-12
+ mcrdlm1d_ca_w_0_140_s_0_840 = 2.91e-05  mcrdlm1d_cc_w_0_140_s_0_840 = 3.59e-11  mcrdlm1d_cf_w_0_140_s_0_840 = 1.16e-11
+ mcrdlm1d_ca_w_0_140_s_1_540 = 2.91e-05  mcrdlm1d_cc_w_0_140_s_1_540 = 2.11e-11  mcrdlm1d_cf_w_0_140_s_1_540 = 1.86e-11
+ mcrdlm1d_ca_w_0_140_s_3_500 = 2.91e-05  mcrdlm1d_cc_w_0_140_s_3_500 = 7.44e-12  mcrdlm1d_cf_w_0_140_s_3_500 = 2.89e-11
+ mcrdlm1d_ca_w_1_120_s_0_140 = 2.91e-05  mcrdlm1d_cc_w_1_120_s_0_140 = 1.12e-10  mcrdlm1d_cf_w_1_120_s_0_140 = 2.50e-12
+ mcrdlm1d_ca_w_1_120_s_0_175 = 2.91e-05  mcrdlm1d_cc_w_1_120_s_0_175 = 1.09e-10  mcrdlm1d_cf_w_1_120_s_0_175 = 3.01e-12
+ mcrdlm1d_ca_w_1_120_s_0_210 = 2.91e-05  mcrdlm1d_cc_w_1_120_s_0_210 = 1.05e-10  mcrdlm1d_cf_w_1_120_s_0_210 = 3.51e-12
+ mcrdlm1d_ca_w_1_120_s_0_280 = 2.91e-05  mcrdlm1d_cc_w_1_120_s_0_280 = 9.31e-11  mcrdlm1d_cf_w_1_120_s_0_280 = 4.51e-12
+ mcrdlm1d_ca_w_1_120_s_0_350 = 2.91e-05  mcrdlm1d_cc_w_1_120_s_0_350 = 8.34e-11  mcrdlm1d_cf_w_1_120_s_0_350 = 5.48e-12
+ mcrdlm1d_ca_w_1_120_s_0_420 = 2.91e-05  mcrdlm1d_cc_w_1_120_s_0_420 = 7.42e-11  mcrdlm1d_cf_w_1_120_s_0_420 = 6.44e-12
+ mcrdlm1d_ca_w_1_120_s_0_560 = 2.91e-05  mcrdlm1d_cc_w_1_120_s_0_560 = 6.17e-11  mcrdlm1d_cf_w_1_120_s_0_560 = 8.29e-12
+ mcrdlm1d_ca_w_1_120_s_0_840 = 2.91e-05  mcrdlm1d_cc_w_1_120_s_0_840 = 4.64e-11  mcrdlm1d_cf_w_1_120_s_0_840 = 1.18e-11
+ mcrdlm1d_ca_w_1_120_s_1_540 = 2.91e-05  mcrdlm1d_cc_w_1_120_s_1_540 = 2.84e-11  mcrdlm1d_cf_w_1_120_s_1_540 = 1.91e-11
+ mcrdlm1d_ca_w_1_120_s_3_500 = 2.91e-05  mcrdlm1d_cc_w_1_120_s_3_500 = 1.10e-11  mcrdlm1d_cf_w_1_120_s_3_500 = 3.11e-11
+ mcrdlm1p1_ca_w_0_140_s_0_140 = 3.48e-05  mcrdlm1p1_cc_w_0_140_s_0_140 = 8.63e-11  mcrdlm1p1_cf_w_0_140_s_0_140 = 2.93e-12
+ mcrdlm1p1_ca_w_0_140_s_0_175 = 3.48e-05  mcrdlm1p1_cc_w_0_140_s_0_175 = 8.47e-11  mcrdlm1p1_cf_w_0_140_s_0_175 = 3.53e-12
+ mcrdlm1p1_ca_w_0_140_s_0_210 = 3.48e-05  mcrdlm1p1_cc_w_0_140_s_0_210 = 8.17e-11  mcrdlm1p1_cf_w_0_140_s_0_210 = 4.14e-12
+ mcrdlm1p1_ca_w_0_140_s_0_280 = 3.48e-05  mcrdlm1p1_cc_w_0_140_s_0_280 = 7.38e-11  mcrdlm1p1_cf_w_0_140_s_0_280 = 5.32e-12
+ mcrdlm1p1_ca_w_0_140_s_0_350 = 3.48e-05  mcrdlm1p1_cc_w_0_140_s_0_350 = 6.48e-11  mcrdlm1p1_cf_w_0_140_s_0_350 = 6.45e-12
+ mcrdlm1p1_ca_w_0_140_s_0_420 = 3.48e-05  mcrdlm1p1_cc_w_0_140_s_0_420 = 5.72e-11  mcrdlm1p1_cf_w_0_140_s_0_420 = 7.62e-12
+ mcrdlm1p1_ca_w_0_140_s_0_560 = 3.48e-05  mcrdlm1p1_cc_w_0_140_s_0_560 = 4.68e-11  mcrdlm1p1_cf_w_0_140_s_0_560 = 9.75e-12
+ mcrdlm1p1_ca_w_0_140_s_0_840 = 3.48e-05  mcrdlm1p1_cc_w_0_140_s_0_840 = 3.43e-11  mcrdlm1p1_cf_w_0_140_s_0_840 = 1.37e-11
+ mcrdlm1p1_ca_w_0_140_s_1_540 = 3.48e-05  mcrdlm1p1_cc_w_0_140_s_1_540 = 1.95e-11  mcrdlm1p1_cf_w_0_140_s_1_540 = 2.14e-11
+ mcrdlm1p1_ca_w_0_140_s_3_500 = 3.48e-05  mcrdlm1p1_cc_w_0_140_s_3_500 = 6.38e-12  mcrdlm1p1_cf_w_0_140_s_3_500 = 3.19e-11
+ mcrdlm1p1_ca_w_1_120_s_0_140 = 3.48e-05  mcrdlm1p1_cc_w_1_120_s_0_140 = 1.10e-10  mcrdlm1p1_cf_w_1_120_s_0_140 = 3.03e-12
+ mcrdlm1p1_ca_w_1_120_s_0_175 = 3.48e-05  mcrdlm1p1_cc_w_1_120_s_0_175 = 1.07e-10  mcrdlm1p1_cf_w_1_120_s_0_175 = 3.64e-12
+ mcrdlm1p1_ca_w_1_120_s_0_210 = 3.48e-05  mcrdlm1p1_cc_w_1_120_s_0_210 = 1.03e-10  mcrdlm1p1_cf_w_1_120_s_0_210 = 4.23e-12
+ mcrdlm1p1_ca_w_1_120_s_0_280 = 3.48e-05  mcrdlm1p1_cc_w_1_120_s_0_280 = 9.10e-11  mcrdlm1p1_cf_w_1_120_s_0_280 = 5.41e-12
+ mcrdlm1p1_ca_w_1_120_s_0_350 = 3.48e-05  mcrdlm1p1_cc_w_1_120_s_0_350 = 8.12e-11  mcrdlm1p1_cf_w_1_120_s_0_350 = 6.57e-12
+ mcrdlm1p1_ca_w_1_120_s_0_420 = 3.48e-05  mcrdlm1p1_cc_w_1_120_s_0_420 = 7.24e-11  mcrdlm1p1_cf_w_1_120_s_0_420 = 7.70e-12
+ mcrdlm1p1_ca_w_1_120_s_0_560 = 3.48e-05  mcrdlm1p1_cc_w_1_120_s_0_560 = 5.95e-11  mcrdlm1p1_cf_w_1_120_s_0_560 = 9.85e-12
+ mcrdlm1p1_ca_w_1_120_s_0_840 = 3.48e-05  mcrdlm1p1_cc_w_1_120_s_0_840 = 4.44e-11  mcrdlm1p1_cf_w_1_120_s_0_840 = 1.39e-11
+ mcrdlm1p1_ca_w_1_120_s_1_540 = 3.48e-05  mcrdlm1p1_cc_w_1_120_s_1_540 = 2.64e-11  mcrdlm1p1_cf_w_1_120_s_1_540 = 2.21e-11
+ mcrdlm1p1_ca_w_1_120_s_3_500 = 3.48e-05  mcrdlm1p1_cc_w_1_120_s_3_500 = 9.76e-12  mcrdlm1p1_cf_w_1_120_s_3_500 = 3.44e-11
+ mcrdlm1l1_ca_w_0_140_s_0_140 = 7.97e-05  mcrdlm1l1_cc_w_0_140_s_0_140 = 8.18e-11  mcrdlm1l1_cf_w_0_140_s_0_140 = 6.43e-12
+ mcrdlm1l1_ca_w_0_140_s_0_175 = 7.97e-05  mcrdlm1l1_cc_w_0_140_s_0_175 = 8.00e-11  mcrdlm1l1_cf_w_0_140_s_0_175 = 7.83e-12
+ mcrdlm1l1_ca_w_0_140_s_0_210 = 7.97e-05  mcrdlm1l1_cc_w_0_140_s_0_210 = 7.65e-11  mcrdlm1l1_cf_w_0_140_s_0_210 = 9.17e-12
+ mcrdlm1l1_ca_w_0_140_s_0_280 = 7.97e-05  mcrdlm1l1_cc_w_0_140_s_0_280 = 6.75e-11  mcrdlm1l1_cf_w_0_140_s_0_280 = 1.17e-11
+ mcrdlm1l1_ca_w_0_140_s_0_350 = 7.97e-05  mcrdlm1l1_cc_w_0_140_s_0_350 = 5.81e-11  mcrdlm1l1_cf_w_0_140_s_0_350 = 1.41e-11
+ mcrdlm1l1_ca_w_0_140_s_0_420 = 7.97e-05  mcrdlm1l1_cc_w_0_140_s_0_420 = 5.04e-11  mcrdlm1l1_cf_w_0_140_s_0_420 = 1.64e-11
+ mcrdlm1l1_ca_w_0_140_s_0_560 = 7.97e-05  mcrdlm1l1_cc_w_0_140_s_0_560 = 3.91e-11  mcrdlm1l1_cf_w_0_140_s_0_560 = 2.06e-11
+ mcrdlm1l1_ca_w_0_140_s_0_840 = 7.97e-05  mcrdlm1l1_cc_w_0_140_s_0_840 = 2.64e-11  mcrdlm1l1_cf_w_0_140_s_0_840 = 2.74e-11
+ mcrdlm1l1_ca_w_0_140_s_1_540 = 7.97e-05  mcrdlm1l1_cc_w_0_140_s_1_540 = 1.24e-11  mcrdlm1l1_cf_w_0_140_s_1_540 = 3.78e-11
+ mcrdlm1l1_ca_w_0_140_s_3_500 = 7.97e-05  mcrdlm1l1_cc_w_0_140_s_3_500 = 3.22e-12  mcrdlm1l1_cf_w_0_140_s_3_500 = 4.66e-11
+ mcrdlm1l1_ca_w_1_120_s_0_140 = 7.97e-05  mcrdlm1l1_cc_w_1_120_s_0_140 = 1.01e-10  mcrdlm1l1_cf_w_1_120_s_0_140 = 6.53e-12
+ mcrdlm1l1_ca_w_1_120_s_0_175 = 7.97e-05  mcrdlm1l1_cc_w_1_120_s_0_175 = 9.75e-11  mcrdlm1l1_cf_w_1_120_s_0_175 = 7.91e-12
+ mcrdlm1l1_ca_w_1_120_s_0_210 = 7.97e-05  mcrdlm1l1_cc_w_1_120_s_0_210 = 9.26e-11  mcrdlm1l1_cf_w_1_120_s_0_210 = 9.24e-12
+ mcrdlm1l1_ca_w_1_120_s_0_280 = 7.97e-05  mcrdlm1l1_cc_w_1_120_s_0_280 = 8.17e-11  mcrdlm1l1_cf_w_1_120_s_0_280 = 1.18e-11
+ mcrdlm1l1_ca_w_1_120_s_0_350 = 7.97e-05  mcrdlm1l1_cc_w_1_120_s_0_350 = 7.15e-11  mcrdlm1l1_cf_w_1_120_s_0_350 = 1.42e-11
+ mcrdlm1l1_ca_w_1_120_s_0_420 = 7.97e-05  mcrdlm1l1_cc_w_1_120_s_0_420 = 6.27e-11  mcrdlm1l1_cf_w_1_120_s_0_420 = 1.65e-11
+ mcrdlm1l1_ca_w_1_120_s_0_560 = 7.97e-05  mcrdlm1l1_cc_w_1_120_s_0_560 = 5.00e-11  mcrdlm1l1_cf_w_1_120_s_0_560 = 2.07e-11
+ mcrdlm1l1_ca_w_1_120_s_0_840 = 7.97e-05  mcrdlm1l1_cc_w_1_120_s_0_840 = 3.52e-11  mcrdlm1l1_cf_w_1_120_s_0_840 = 2.76e-11
+ mcrdlm1l1_ca_w_1_120_s_1_540 = 7.97e-05  mcrdlm1l1_cc_w_1_120_s_1_540 = 1.87e-11  mcrdlm1l1_cf_w_1_120_s_1_540 = 3.89e-11
+ mcrdlm1l1_ca_w_1_120_s_3_500 = 7.97e-05  mcrdlm1l1_cc_w_1_120_s_3_500 = 5.85e-12  mcrdlm1l1_cf_w_1_120_s_3_500 = 5.05e-11
+ mcm3m2f_ca_w_0_140_s_0_140 = 7.34e-05  mcm3m2f_cc_w_0_140_s_0_140 = 8.24e-11  mcm3m2f_cf_w_0_140_s_0_140 = 5.92e-12
+ mcm3m2f_ca_w_0_140_s_0_175 = 7.34e-05  mcm3m2f_cc_w_0_140_s_0_175 = 8.11e-11  mcm3m2f_cf_w_0_140_s_0_175 = 7.08e-12
+ mcm3m2f_ca_w_0_140_s_0_210 = 7.34e-05  mcm3m2f_cc_w_0_140_s_0_210 = 7.70e-11  mcm3m2f_cf_w_0_140_s_0_210 = 8.28e-12
+ mcm3m2f_ca_w_0_140_s_0_280 = 7.34e-05  mcm3m2f_cc_w_0_140_s_0_280 = 6.80e-11  mcm3m2f_cf_w_0_140_s_0_280 = 1.05e-11
+ mcm3m2f_ca_w_0_140_s_0_350 = 7.34e-05  mcm3m2f_cc_w_0_140_s_0_350 = 5.84e-11  mcm3m2f_cf_w_0_140_s_0_350 = 1.27e-11
+ mcm3m2f_ca_w_0_140_s_0_420 = 7.34e-05  mcm3m2f_cc_w_0_140_s_0_420 = 5.06e-11  mcm3m2f_cf_w_0_140_s_0_420 = 1.48e-11
+ mcm3m2f_ca_w_0_140_s_0_560 = 7.34e-05  mcm3m2f_cc_w_0_140_s_0_560 = 3.91e-11  mcm3m2f_cf_w_0_140_s_0_560 = 1.87e-11
+ mcm3m2f_ca_w_0_140_s_0_840 = 7.34e-05  mcm3m2f_cc_w_0_140_s_0_840 = 2.55e-11  mcm3m2f_cf_w_0_140_s_0_840 = 2.52e-11
+ mcm3m2f_ca_w_0_140_s_1_540 = 7.34e-05  mcm3m2f_cc_w_0_140_s_1_540 = 1.05e-11  mcm3m2f_cf_w_0_140_s_1_540 = 3.55e-11
+ mcm3m2f_ca_w_0_140_s_3_500 = 7.34e-05  mcm3m2f_cc_w_0_140_s_3_500 = 1.43e-12  mcm3m2f_cf_w_0_140_s_3_500 = 4.37e-11
+ mcm3m2f_ca_w_1_120_s_0_140 = 7.34e-05  mcm3m2f_cc_w_1_120_s_0_140 = 9.69e-11  mcm3m2f_cf_w_1_120_s_0_140 = 5.96e-12
+ mcm3m2f_ca_w_1_120_s_0_175 = 7.34e-05  mcm3m2f_cc_w_1_120_s_0_175 = 9.45e-11  mcm3m2f_cf_w_1_120_s_0_175 = 7.13e-12
+ mcm3m2f_ca_w_1_120_s_0_210 = 7.34e-05  mcm3m2f_cc_w_1_120_s_0_210 = 8.96e-11  mcm3m2f_cf_w_1_120_s_0_210 = 8.29e-12
+ mcm3m2f_ca_w_1_120_s_0_280 = 7.34e-05  mcm3m2f_cc_w_1_120_s_0_280 = 7.87e-11  mcm3m2f_cf_w_1_120_s_0_280 = 1.06e-11
+ mcm3m2f_ca_w_1_120_s_0_350 = 7.34e-05  mcm3m2f_cc_w_1_120_s_0_350 = 6.79e-11  mcm3m2f_cf_w_1_120_s_0_350 = 1.28e-11
+ mcm3m2f_ca_w_1_120_s_0_420 = 7.34e-05  mcm3m2f_cc_w_1_120_s_0_420 = 5.88e-11  mcm3m2f_cf_w_1_120_s_0_420 = 1.49e-11
+ mcm3m2f_ca_w_1_120_s_0_560 = 7.34e-05  mcm3m2f_cc_w_1_120_s_0_560 = 4.57e-11  mcm3m2f_cf_w_1_120_s_0_560 = 1.89e-11
+ mcm3m2f_ca_w_1_120_s_0_840 = 7.34e-05  mcm3m2f_cc_w_1_120_s_0_840 = 3.01e-11  mcm3m2f_cf_w_1_120_s_0_840 = 2.56e-11
+ mcm3m2f_ca_w_1_120_s_1_540 = 7.34e-05  mcm3m2f_cc_w_1_120_s_1_540 = 1.31e-11  mcm3m2f_cf_w_1_120_s_1_540 = 3.68e-11
+ mcm3m2f_ca_w_1_120_s_3_500 = 7.34e-05  mcm3m2f_cc_w_1_120_s_3_500 = 1.89e-12  mcm3m2f_cf_w_1_120_s_3_500 = 4.67e-11
+ mcm3m2d_ca_w_0_140_s_0_140 = 7.63e-05  mcm3m2d_cc_w_0_140_s_0_140 = 8.21e-11  mcm3m2d_cf_w_0_140_s_0_140 = 6.15e-12
+ mcm3m2d_ca_w_0_140_s_0_175 = 7.63e-05  mcm3m2d_cc_w_0_140_s_0_175 = 8.07e-11  mcm3m2d_cf_w_0_140_s_0_175 = 7.37e-12
+ mcm3m2d_ca_w_0_140_s_0_210 = 7.63e-05  mcm3m2d_cc_w_0_140_s_0_210 = 7.68e-11  mcm3m2d_cf_w_0_140_s_0_210 = 8.62e-12
+ mcm3m2d_ca_w_0_140_s_0_280 = 7.63e-05  mcm3m2d_cc_w_0_140_s_0_280 = 6.75e-11  mcm3m2d_cf_w_0_140_s_0_280 = 1.09e-11
+ mcm3m2d_ca_w_0_140_s_0_350 = 7.63e-05  mcm3m2d_cc_w_0_140_s_0_350 = 5.79e-11  mcm3m2d_cf_w_0_140_s_0_350 = 1.32e-11
+ mcm3m2d_ca_w_0_140_s_0_420 = 7.63e-05  mcm3m2d_cc_w_0_140_s_0_420 = 4.98e-11  mcm3m2d_cf_w_0_140_s_0_420 = 1.54e-11
+ mcm3m2d_ca_w_0_140_s_0_560 = 7.63e-05  mcm3m2d_cc_w_0_140_s_0_560 = 3.83e-11  mcm3m2d_cf_w_0_140_s_0_560 = 1.94e-11
+ mcm3m2d_ca_w_0_140_s_0_840 = 7.63e-05  mcm3m2d_cc_w_0_140_s_0_840 = 2.46e-11  mcm3m2d_cf_w_0_140_s_0_840 = 2.61e-11
+ mcm3m2d_ca_w_0_140_s_1_540 = 7.63e-05  mcm3m2d_cc_w_0_140_s_1_540 = 9.65e-12  mcm3m2d_cf_w_0_140_s_1_540 = 3.66e-11
+ mcm3m2d_ca_w_0_140_s_3_500 = 7.63e-05  mcm3m2d_cc_w_0_140_s_3_500 = 1.09e-12  mcm3m2d_cf_w_0_140_s_3_500 = 4.45e-11
+ mcm3m2d_ca_w_1_120_s_0_140 = 7.63e-05  mcm3m2d_cc_w_1_120_s_0_140 = 9.58e-11  mcm3m2d_cf_w_1_120_s_0_140 = 6.20e-12
+ mcm3m2d_ca_w_1_120_s_0_175 = 7.63e-05  mcm3m2d_cc_w_1_120_s_0_175 = 9.32e-11  mcm3m2d_cf_w_1_120_s_0_175 = 7.42e-12
+ mcm3m2d_ca_w_1_120_s_0_210 = 7.63e-05  mcm3m2d_cc_w_1_120_s_0_210 = 8.84e-11  mcm3m2d_cf_w_1_120_s_0_210 = 8.63e-12
+ mcm3m2d_ca_w_1_120_s_0_280 = 7.63e-05  mcm3m2d_cc_w_1_120_s_0_280 = 7.73e-11  mcm3m2d_cf_w_1_120_s_0_280 = 1.10e-11
+ mcm3m2d_ca_w_1_120_s_0_350 = 7.63e-05  mcm3m2d_cc_w_1_120_s_0_350 = 6.64e-11  mcm3m2d_cf_w_1_120_s_0_350 = 1.33e-11
+ mcm3m2d_ca_w_1_120_s_0_420 = 7.63e-05  mcm3m2d_cc_w_1_120_s_0_420 = 5.73e-11  mcm3m2d_cf_w_1_120_s_0_420 = 1.56e-11
+ mcm3m2d_ca_w_1_120_s_0_560 = 7.63e-05  mcm3m2d_cc_w_1_120_s_0_560 = 4.42e-11  mcm3m2d_cf_w_1_120_s_0_560 = 1.96e-11
+ mcm3m2d_ca_w_1_120_s_0_840 = 7.63e-05  mcm3m2d_cc_w_1_120_s_0_840 = 2.86e-11  mcm3m2d_cf_w_1_120_s_0_840 = 2.66e-11
+ mcm3m2d_ca_w_1_120_s_1_540 = 7.63e-05  mcm3m2d_cc_w_1_120_s_1_540 = 1.17e-11  mcm3m2d_cf_w_1_120_s_1_540 = 3.79e-11
+ mcm3m2d_ca_w_1_120_s_3_500 = 7.63e-05  mcm3m2d_cc_w_1_120_s_3_500 = 1.42e-12  mcm3m2d_cf_w_1_120_s_3_500 = 4.72e-11
+ mcm3m2p1_ca_w_0_140_s_0_140 = 7.84e-05  mcm3m2p1_cc_w_0_140_s_0_140 = 8.19e-11  mcm3m2p1_cf_w_0_140_s_0_140 = 6.33e-12
+ mcm3m2p1_ca_w_0_140_s_0_175 = 7.84e-05  mcm3m2p1_cc_w_0_140_s_0_175 = 8.01e-11  mcm3m2p1_cf_w_0_140_s_0_175 = 7.59e-12
+ mcm3m2p1_ca_w_0_140_s_0_210 = 7.84e-05  mcm3m2p1_cc_w_0_140_s_0_210 = 7.63e-11  mcm3m2p1_cf_w_0_140_s_0_210 = 8.85e-12
+ mcm3m2p1_ca_w_0_140_s_0_280 = 7.84e-05  mcm3m2p1_cc_w_0_140_s_0_280 = 6.71e-11  mcm3m2p1_cf_w_0_140_s_0_280 = 1.12e-11
+ mcm3m2p1_ca_w_0_140_s_0_350 = 7.84e-05  mcm3m2p1_cc_w_0_140_s_0_350 = 5.75e-11  mcm3m2p1_cf_w_0_140_s_0_350 = 1.36e-11
+ mcm3m2p1_ca_w_0_140_s_0_420 = 7.84e-05  mcm3m2p1_cc_w_0_140_s_0_420 = 4.94e-11  mcm3m2p1_cf_w_0_140_s_0_420 = 1.59e-11
+ mcm3m2p1_ca_w_0_140_s_0_560 = 7.84e-05  mcm3m2p1_cc_w_0_140_s_0_560 = 3.78e-11  mcm3m2p1_cf_w_0_140_s_0_560 = 1.99e-11
+ mcm3m2p1_ca_w_0_140_s_0_840 = 7.84e-05  mcm3m2p1_cc_w_0_140_s_0_840 = 2.39e-11  mcm3m2p1_cf_w_0_140_s_0_840 = 2.68e-11
+ mcm3m2p1_ca_w_0_140_s_1_540 = 7.84e-05  mcm3m2p1_cc_w_0_140_s_1_540 = 9.11e-12  mcm3m2p1_cf_w_0_140_s_1_540 = 3.75e-11
+ mcm3m2p1_ca_w_0_140_s_3_500 = 7.84e-05  mcm3m2p1_cc_w_0_140_s_3_500 = 9.15e-13  mcm3m2p1_cf_w_0_140_s_3_500 = 4.50e-11
+ mcm3m2p1_ca_w_1_120_s_0_140 = 7.84e-05  mcm3m2p1_cc_w_1_120_s_0_140 = 9.53e-11  mcm3m2p1_cf_w_1_120_s_0_140 = 6.39e-12
+ mcm3m2p1_ca_w_1_120_s_0_175 = 7.84e-05  mcm3m2p1_cc_w_1_120_s_0_175 = 9.22e-11  mcm3m2p1_cf_w_1_120_s_0_175 = 7.65e-12
+ mcm3m2p1_ca_w_1_120_s_0_210 = 7.84e-05  mcm3m2p1_cc_w_1_120_s_0_210 = 8.74e-11  mcm3m2p1_cf_w_1_120_s_0_210 = 8.90e-12
+ mcm3m2p1_ca_w_1_120_s_0_280 = 7.84e-05  mcm3m2p1_cc_w_1_120_s_0_280 = 7.62e-11  mcm3m2p1_cf_w_1_120_s_0_280 = 1.13e-11
+ mcm3m2p1_ca_w_1_120_s_0_350 = 7.84e-05  mcm3m2p1_cc_w_1_120_s_0_350 = 6.55e-11  mcm3m2p1_cf_w_1_120_s_0_350 = 1.37e-11
+ mcm3m2p1_ca_w_1_120_s_0_420 = 7.84e-05  mcm3m2p1_cc_w_1_120_s_0_420 = 5.62e-11  mcm3m2p1_cf_w_1_120_s_0_420 = 1.60e-11
+ mcm3m2p1_ca_w_1_120_s_0_560 = 7.84e-05  mcm3m2p1_cc_w_1_120_s_0_560 = 4.31e-11  mcm3m2p1_cf_w_1_120_s_0_560 = 2.02e-11
+ mcm3m2p1_ca_w_1_120_s_0_840 = 7.84e-05  mcm3m2p1_cc_w_1_120_s_0_840 = 2.76e-11  mcm3m2p1_cf_w_1_120_s_0_840 = 2.73e-11
+ mcm3m2p1_ca_w_1_120_s_1_540 = 7.84e-05  mcm3m2p1_cc_w_1_120_s_1_540 = 1.09e-11  mcm3m2p1_cf_w_1_120_s_1_540 = 3.88e-11
+ mcm3m2p1_ca_w_1_120_s_3_500 = 7.84e-05  mcm3m2p1_cc_w_1_120_s_3_500 = 1.08e-12  mcm3m2p1_cf_w_1_120_s_3_500 = 4.76e-11
+ mcm3m2l1_ca_w_0_140_s_0_140 = 8.81e-05  mcm3m2l1_cc_w_0_140_s_0_140 = 8.08e-11  mcm3m2l1_cf_w_0_140_s_0_140 = 7.12e-12
+ mcm3m2l1_ca_w_0_140_s_0_175 = 8.81e-05  mcm3m2l1_cc_w_0_140_s_0_175 = 7.89e-11  mcm3m2l1_cf_w_0_140_s_0_175 = 8.55e-12
+ mcm3m2l1_ca_w_0_140_s_0_210 = 8.81e-05  mcm3m2l1_cc_w_0_140_s_0_210 = 7.50e-11  mcm3m2l1_cf_w_0_140_s_0_210 = 9.97e-12
+ mcm3m2l1_ca_w_0_140_s_0_280 = 8.81e-05  mcm3m2l1_cc_w_0_140_s_0_280 = 6.55e-11  mcm3m2l1_cf_w_0_140_s_0_280 = 1.27e-11
+ mcm3m2l1_ca_w_0_140_s_0_350 = 8.81e-05  mcm3m2l1_cc_w_0_140_s_0_350 = 5.58e-11  mcm3m2l1_cf_w_0_140_s_0_350 = 1.53e-11
+ mcm3m2l1_ca_w_0_140_s_0_420 = 8.81e-05  mcm3m2l1_cc_w_0_140_s_0_420 = 4.71e-11  mcm3m2l1_cf_w_0_140_s_0_420 = 1.79e-11
+ mcm3m2l1_ca_w_0_140_s_0_560 = 8.81e-05  mcm3m2l1_cc_w_0_140_s_0_560 = 3.56e-11  mcm3m2l1_cf_w_0_140_s_0_560 = 2.24e-11
+ mcm3m2l1_ca_w_0_140_s_0_840 = 8.81e-05  mcm3m2l1_cc_w_0_140_s_0_840 = 2.14e-11  mcm3m2l1_cf_w_0_140_s_0_840 = 3.00e-11
+ mcm3m2l1_ca_w_0_140_s_1_540 = 8.81e-05  mcm3m2l1_cc_w_0_140_s_1_540 = 7.00e-12  mcm3m2l1_cf_w_0_140_s_1_540 = 4.09e-11
+ mcm3m2l1_ca_w_0_140_s_3_500 = 8.81e-05  mcm3m2l1_cc_w_0_140_s_3_500 = 4.15e-13  mcm3m2l1_cf_w_0_140_s_3_500 = 4.71e-11
+ mcm3m2l1_ca_w_1_120_s_0_140 = 8.81e-05  mcm3m2l1_cc_w_1_120_s_0_140 = 9.14e-11  mcm3m2l1_cf_w_1_120_s_0_140 = 7.17e-12
+ mcm3m2l1_ca_w_1_120_s_0_175 = 8.81e-05  mcm3m2l1_cc_w_1_120_s_0_175 = 8.88e-11  mcm3m2l1_cf_w_1_120_s_0_175 = 8.60e-12
+ mcm3m2l1_ca_w_1_120_s_0_210 = 8.81e-05  mcm3m2l1_cc_w_1_120_s_0_210 = 8.38e-11  mcm3m2l1_cf_w_1_120_s_0_210 = 1.00e-11
+ mcm3m2l1_ca_w_1_120_s_0_280 = 8.81e-05  mcm3m2l1_cc_w_1_120_s_0_280 = 7.24e-11  mcm3m2l1_cf_w_1_120_s_0_280 = 1.27e-11
+ mcm3m2l1_ca_w_1_120_s_0_350 = 8.81e-05  mcm3m2l1_cc_w_1_120_s_0_350 = 6.17e-11  mcm3m2l1_cf_w_1_120_s_0_350 = 1.54e-11
+ mcm3m2l1_ca_w_1_120_s_0_420 = 8.81e-05  mcm3m2l1_cc_w_1_120_s_0_420 = 5.24e-11  mcm3m2l1_cf_w_1_120_s_0_420 = 1.81e-11
+ mcm3m2l1_ca_w_1_120_s_0_560 = 8.81e-05  mcm3m2l1_cc_w_1_120_s_0_560 = 3.91e-11  mcm3m2l1_cf_w_1_120_s_0_560 = 2.27e-11
+ mcm3m2l1_ca_w_1_120_s_0_840 = 8.81e-05  mcm3m2l1_cc_w_1_120_s_0_840 = 2.37e-11  mcm3m2l1_cf_w_1_120_s_0_840 = 3.05e-11
+ mcm3m2l1_ca_w_1_120_s_1_540 = 8.81e-05  mcm3m2l1_cc_w_1_120_s_1_540 = 7.86e-12  mcm3m2l1_cf_w_1_120_s_1_540 = 4.21e-11
+ mcm3m2l1_ca_w_1_120_s_3_500 = 8.81e-05  mcm3m2l1_cc_w_1_120_s_3_500 = 4.95e-13  mcm3m2l1_cf_w_1_120_s_3_500 = 4.92e-11
+ mcm3m2m1_ca_w_0_140_s_0_140 = 1.40e-04  mcm3m2m1_cc_w_0_140_s_0_140 = 7.47e-11  mcm3m2m1_cf_w_0_140_s_0_140 = 1.12e-11
+ mcm3m2m1_ca_w_0_140_s_0_175 = 1.40e-04  mcm3m2m1_cc_w_0_140_s_0_175 = 7.33e-11  mcm3m2m1_cf_w_0_140_s_0_175 = 1.35e-11
+ mcm3m2m1_ca_w_0_140_s_0_210 = 1.40e-04  mcm3m2m1_cc_w_0_140_s_0_210 = 6.89e-11  mcm3m2m1_cf_w_0_140_s_0_210 = 1.57e-11
+ mcm3m2m1_ca_w_0_140_s_0_280 = 1.40e-04  mcm3m2m1_cc_w_0_140_s_0_280 = 5.86e-11  mcm3m2m1_cf_w_0_140_s_0_280 = 2.00e-11
+ mcm3m2m1_ca_w_0_140_s_0_350 = 1.40e-04  mcm3m2m1_cc_w_0_140_s_0_350 = 4.82e-11  mcm3m2m1_cf_w_0_140_s_0_350 = 2.42e-11
+ mcm3m2m1_ca_w_0_140_s_0_420 = 1.40e-04  mcm3m2m1_cc_w_0_140_s_0_420 = 3.96e-11  mcm3m2m1_cf_w_0_140_s_0_420 = 2.78e-11
+ mcm3m2m1_ca_w_0_140_s_0_560 = 1.40e-04  mcm3m2m1_cc_w_0_140_s_0_560 = 2.73e-11  mcm3m2m1_cf_w_0_140_s_0_560 = 3.44e-11
+ mcm3m2m1_ca_w_0_140_s_0_840 = 1.40e-04  mcm3m2m1_cc_w_0_140_s_0_840 = 1.37e-11  mcm3m2m1_cf_w_0_140_s_0_840 = 4.39e-11
+ mcm3m2m1_ca_w_0_140_s_1_540 = 1.40e-04  mcm3m2m1_cc_w_0_140_s_1_540 = 2.64e-12  mcm3m2m1_cf_w_0_140_s_1_540 = 5.40e-11
+ mcm3m2m1_ca_w_0_140_s_3_500 = 1.40e-04  mcm3m2m1_cc_w_0_140_s_3_500 = 6.00e-14  mcm3m2m1_cf_w_0_140_s_3_500 = 5.72e-11
+ mcm3m2m1_ca_w_1_120_s_0_140 = 1.40e-04  mcm3m2m1_cc_w_1_120_s_0_140 = 8.02e-11  mcm3m2m1_cf_w_1_120_s_0_140 = 1.12e-11
+ mcm3m2m1_ca_w_1_120_s_0_175 = 1.40e-04  mcm3m2m1_cc_w_1_120_s_0_175 = 7.77e-11  mcm3m2m1_cf_w_1_120_s_0_175 = 1.35e-11
+ mcm3m2m1_ca_w_1_120_s_0_210 = 1.40e-04  mcm3m2m1_cc_w_1_120_s_0_210 = 7.30e-11  mcm3m2m1_cf_w_1_120_s_0_210 = 1.58e-11
+ mcm3m2m1_ca_w_1_120_s_0_280 = 1.40e-04  mcm3m2m1_cc_w_1_120_s_0_280 = 6.13e-11  mcm3m2m1_cf_w_1_120_s_0_280 = 2.01e-11
+ mcm3m2m1_ca_w_1_120_s_0_350 = 1.40e-04  mcm3m2m1_cc_w_1_120_s_0_350 = 5.07e-11  mcm3m2m1_cf_w_1_120_s_0_350 = 2.42e-11
+ mcm3m2m1_ca_w_1_120_s_0_420 = 1.40e-04  mcm3m2m1_cc_w_1_120_s_0_420 = 4.17e-11  mcm3m2m1_cf_w_1_120_s_0_420 = 2.81e-11
+ mcm3m2m1_ca_w_1_120_s_0_560 = 1.40e-04  mcm3m2m1_cc_w_1_120_s_0_560 = 2.89e-11  mcm3m2m1_cf_w_1_120_s_0_560 = 3.47e-11
+ mcm3m2m1_ca_w_1_120_s_0_840 = 1.40e-04  mcm3m2m1_cc_w_1_120_s_0_840 = 1.44e-11  mcm3m2m1_cf_w_1_120_s_0_840 = 4.45e-11
+ mcm3m2m1_ca_w_1_120_s_1_540 = 1.40e-04  mcm3m2m1_cc_w_1_120_s_1_540 = 2.85e-12  mcm3m2m1_cf_w_1_120_s_1_540 = 5.51e-11
+ mcm3m2m1_ca_w_1_120_s_3_500 = 1.40e-04  mcm3m2m1_cc_w_1_120_s_3_500 = 1.00e-13  mcm3m2m1_cf_w_1_120_s_3_500 = 5.82e-11
+ mcm4m2f_ca_w_0_140_s_0_140 = 3.17e-05  mcm4m2f_cc_w_0_140_s_0_140 = 8.69e-11  mcm4m2f_cf_w_0_140_s_0_140 = 2.67e-12
+ mcm4m2f_ca_w_0_140_s_0_175 = 3.17e-05  mcm4m2f_cc_w_0_140_s_0_175 = 8.55e-11  mcm4m2f_cf_w_0_140_s_0_175 = 3.21e-12
+ mcm4m2f_ca_w_0_140_s_0_210 = 3.17e-05  mcm4m2f_cc_w_0_140_s_0_210 = 8.23e-11  mcm4m2f_cf_w_0_140_s_0_210 = 3.79e-12
+ mcm4m2f_ca_w_0_140_s_0_280 = 3.17e-05  mcm4m2f_cc_w_0_140_s_0_280 = 7.42e-11  mcm4m2f_cf_w_0_140_s_0_280 = 4.84e-12
+ mcm4m2f_ca_w_0_140_s_0_350 = 3.17e-05  mcm4m2f_cc_w_0_140_s_0_350 = 6.52e-11  mcm4m2f_cf_w_0_140_s_0_350 = 5.89e-12
+ mcm4m2f_ca_w_0_140_s_0_420 = 3.17e-05  mcm4m2f_cc_w_0_140_s_0_420 = 5.78e-11  mcm4m2f_cf_w_0_140_s_0_420 = 6.98e-12
+ mcm4m2f_ca_w_0_140_s_0_560 = 3.17e-05  mcm4m2f_cc_w_0_140_s_0_560 = 4.72e-11  mcm4m2f_cf_w_0_140_s_0_560 = 8.99e-12
+ mcm4m2f_ca_w_0_140_s_0_840 = 3.17e-05  mcm4m2f_cc_w_0_140_s_0_840 = 3.43e-11  mcm4m2f_cf_w_0_140_s_0_840 = 1.27e-11
+ mcm4m2f_ca_w_0_140_s_1_540 = 3.17e-05  mcm4m2f_cc_w_0_140_s_1_540 = 1.85e-11  mcm4m2f_cf_w_0_140_s_1_540 = 2.02e-11
+ mcm4m2f_ca_w_0_140_s_3_500 = 3.17e-05  mcm4m2f_cc_w_0_140_s_3_500 = 4.59e-12  mcm4m2f_cf_w_0_140_s_3_500 = 3.06e-11
+ mcm4m2f_ca_w_1_120_s_0_140 = 3.17e-05  mcm4m2f_cc_w_1_120_s_0_140 = 1.09e-10  mcm4m2f_cf_w_1_120_s_0_140 = 2.69e-12
+ mcm4m2f_ca_w_1_120_s_0_175 = 3.17e-05  mcm4m2f_cc_w_1_120_s_0_175 = 1.06e-10  mcm4m2f_cf_w_1_120_s_0_175 = 3.24e-12
+ mcm4m2f_ca_w_1_120_s_0_210 = 3.17e-05  mcm4m2f_cc_w_1_120_s_0_210 = 1.02e-10  mcm4m2f_cf_w_1_120_s_0_210 = 3.78e-12
+ mcm4m2f_ca_w_1_120_s_0_280 = 3.17e-05  mcm4m2f_cc_w_1_120_s_0_280 = 9.03e-11  mcm4m2f_cf_w_1_120_s_0_280 = 4.87e-12
+ mcm4m2f_ca_w_1_120_s_0_350 = 3.17e-05  mcm4m2f_cc_w_1_120_s_0_350 = 7.97e-11  mcm4m2f_cf_w_1_120_s_0_350 = 5.92e-12
+ mcm4m2f_ca_w_1_120_s_0_420 = 3.17e-05  mcm4m2f_cc_w_1_120_s_0_420 = 7.09e-11  mcm4m2f_cf_w_1_120_s_0_420 = 6.99e-12
+ mcm4m2f_ca_w_1_120_s_0_560 = 3.17e-05  mcm4m2f_cc_w_1_120_s_0_560 = 5.78e-11  mcm4m2f_cf_w_1_120_s_0_560 = 9.00e-12
+ mcm4m2f_ca_w_1_120_s_0_840 = 3.17e-05  mcm4m2f_cc_w_1_120_s_0_840 = 4.18e-11  mcm4m2f_cf_w_1_120_s_0_840 = 1.28e-11
+ mcm4m2f_ca_w_1_120_s_1_540 = 3.17e-05  mcm4m2f_cc_w_1_120_s_1_540 = 2.29e-11  mcm4m2f_cf_w_1_120_s_1_540 = 2.09e-11
+ mcm4m2f_ca_w_1_120_s_3_500 = 3.17e-05  mcm4m2f_cc_w_1_120_s_3_500 = 5.85e-12  mcm4m2f_cf_w_1_120_s_3_500 = 3.30e-11
+ mcm4m2d_ca_w_0_140_s_0_140 = 3.46e-05  mcm4m2d_cc_w_0_140_s_0_140 = 8.62e-11  mcm4m2d_cf_w_0_140_s_0_140 = 2.91e-12
+ mcm4m2d_ca_w_0_140_s_0_175 = 3.46e-05  mcm4m2d_cc_w_0_140_s_0_175 = 8.51e-11  mcm4m2d_cf_w_0_140_s_0_175 = 3.49e-12
+ mcm4m2d_ca_w_0_140_s_0_210 = 3.46e-05  mcm4m2d_cc_w_0_140_s_0_210 = 8.19e-11  mcm4m2d_cf_w_0_140_s_0_210 = 4.13e-12
+ mcm4m2d_ca_w_0_140_s_0_280 = 3.46e-05  mcm4m2d_cc_w_0_140_s_0_280 = 7.38e-11  mcm4m2d_cf_w_0_140_s_0_280 = 5.27e-12
+ mcm4m2d_ca_w_0_140_s_0_350 = 3.46e-05  mcm4m2d_cc_w_0_140_s_0_350 = 6.47e-11  mcm4m2d_cf_w_0_140_s_0_350 = 6.41e-12
+ mcm4m2d_ca_w_0_140_s_0_420 = 3.46e-05  mcm4m2d_cc_w_0_140_s_0_420 = 5.72e-11  mcm4m2d_cf_w_0_140_s_0_420 = 7.59e-12
+ mcm4m2d_ca_w_0_140_s_0_560 = 3.46e-05  mcm4m2d_cc_w_0_140_s_0_560 = 4.64e-11  mcm4m2d_cf_w_0_140_s_0_560 = 9.77e-12
+ mcm4m2d_ca_w_0_140_s_0_840 = 3.46e-05  mcm4m2d_cc_w_0_140_s_0_840 = 3.32e-11  mcm4m2d_cf_w_0_140_s_0_840 = 1.37e-11
+ mcm4m2d_ca_w_0_140_s_1_540 = 3.46e-05  mcm4m2d_cc_w_0_140_s_1_540 = 1.74e-11  mcm4m2d_cf_w_0_140_s_1_540 = 2.17e-11
+ mcm4m2d_ca_w_0_140_s_3_500 = 3.46e-05  mcm4m2d_cc_w_0_140_s_3_500 = 3.88e-12  mcm4m2d_cf_w_0_140_s_3_500 = 3.20e-11
+ mcm4m2d_ca_w_1_120_s_0_140 = 3.46e-05  mcm4m2d_cc_w_1_120_s_0_140 = 1.08e-10  mcm4m2d_cf_w_1_120_s_0_140 = 2.93e-12
+ mcm4m2d_ca_w_1_120_s_0_175 = 3.46e-05  mcm4m2d_cc_w_1_120_s_0_175 = 1.05e-10  mcm4m2d_cf_w_1_120_s_0_175 = 3.53e-12
+ mcm4m2d_ca_w_1_120_s_0_210 = 3.46e-05  mcm4m2d_cc_w_1_120_s_0_210 = 1.01e-10  mcm4m2d_cf_w_1_120_s_0_210 = 4.12e-12
+ mcm4m2d_ca_w_1_120_s_0_280 = 3.46e-05  mcm4m2d_cc_w_1_120_s_0_280 = 8.95e-11  mcm4m2d_cf_w_1_120_s_0_280 = 5.29e-12
+ mcm4m2d_ca_w_1_120_s_0_350 = 3.46e-05  mcm4m2d_cc_w_1_120_s_0_350 = 7.84e-11  mcm4m2d_cf_w_1_120_s_0_350 = 6.45e-12
+ mcm4m2d_ca_w_1_120_s_0_420 = 3.46e-05  mcm4m2d_cc_w_1_120_s_0_420 = 6.95e-11  mcm4m2d_cf_w_1_120_s_0_420 = 7.61e-12
+ mcm4m2d_ca_w_1_120_s_0_560 = 3.46e-05  mcm4m2d_cc_w_1_120_s_0_560 = 5.62e-11  mcm4m2d_cf_w_1_120_s_0_560 = 9.79e-12
+ mcm4m2d_ca_w_1_120_s_0_840 = 3.46e-05  mcm4m2d_cc_w_1_120_s_0_840 = 4.02e-11  mcm4m2d_cf_w_1_120_s_0_840 = 1.39e-11
+ mcm4m2d_ca_w_1_120_s_1_540 = 3.46e-05  mcm4m2d_cc_w_1_120_s_1_540 = 2.13e-11  mcm4m2d_cf_w_1_120_s_1_540 = 2.24e-11
+ mcm4m2d_ca_w_1_120_s_3_500 = 3.46e-05  mcm4m2d_cc_w_1_120_s_3_500 = 4.88e-12  mcm4m2d_cf_w_1_120_s_3_500 = 3.45e-11
+ mcm4m2p1_ca_w_0_140_s_0_140 = 3.67e-05  mcm4m2p1_cc_w_0_140_s_0_140 = 8.62e-11  mcm4m2p1_cf_w_0_140_s_0_140 = 3.09e-12
+ mcm4m2p1_ca_w_0_140_s_0_175 = 3.67e-05  mcm4m2p1_cc_w_0_140_s_0_175 = 8.49e-11  mcm4m2p1_cf_w_0_140_s_0_175 = 3.71e-12
+ mcm4m2p1_ca_w_0_140_s_0_210 = 3.67e-05  mcm4m2p1_cc_w_0_140_s_0_210 = 8.14e-11  mcm4m2p1_cf_w_0_140_s_0_210 = 4.38e-12
+ mcm4m2p1_ca_w_0_140_s_0_280 = 3.67e-05  mcm4m2p1_cc_w_0_140_s_0_280 = 7.34e-11  mcm4m2p1_cf_w_0_140_s_0_280 = 5.59e-12
+ mcm4m2p1_ca_w_0_140_s_0_350 = 3.67e-05  mcm4m2p1_cc_w_0_140_s_0_350 = 6.44e-11  mcm4m2p1_cf_w_0_140_s_0_350 = 6.80e-12
+ mcm4m2p1_ca_w_0_140_s_0_420 = 3.67e-05  mcm4m2p1_cc_w_0_140_s_0_420 = 5.65e-11  mcm4m2p1_cf_w_0_140_s_0_420 = 8.05e-12
+ mcm4m2p1_ca_w_0_140_s_0_560 = 3.67e-05  mcm4m2p1_cc_w_0_140_s_0_560 = 4.57e-11  mcm4m2p1_cf_w_0_140_s_0_560 = 1.03e-11
+ mcm4m2p1_ca_w_0_140_s_0_840 = 3.67e-05  mcm4m2p1_cc_w_0_140_s_0_840 = 3.26e-11  mcm4m2p1_cf_w_0_140_s_0_840 = 1.45e-11
+ mcm4m2p1_ca_w_0_140_s_1_540 = 3.67e-05  mcm4m2p1_cc_w_0_140_s_1_540 = 1.66e-11  mcm4m2p1_cf_w_0_140_s_1_540 = 2.27e-11
+ mcm4m2p1_ca_w_0_140_s_3_500 = 3.67e-05  mcm4m2p1_cc_w_0_140_s_3_500 = 3.45e-12  mcm4m2p1_cf_w_0_140_s_3_500 = 3.31e-11
+ mcm4m2p1_ca_w_1_120_s_0_140 = 3.67e-05  mcm4m2p1_cc_w_1_120_s_0_140 = 1.07e-10  mcm4m2p1_cf_w_1_120_s_0_140 = 3.13e-12
+ mcm4m2p1_ca_w_1_120_s_0_175 = 3.67e-05  mcm4m2p1_cc_w_1_120_s_0_175 = 1.04e-10  mcm4m2p1_cf_w_1_120_s_0_175 = 3.76e-12
+ mcm4m2p1_ca_w_1_120_s_0_210 = 3.67e-05  mcm4m2p1_cc_w_1_120_s_0_210 = 9.92e-11  mcm4m2p1_cf_w_1_120_s_0_210 = 4.39e-12
+ mcm4m2p1_ca_w_1_120_s_0_280 = 3.67e-05  mcm4m2p1_cc_w_1_120_s_0_280 = 8.80e-11  mcm4m2p1_cf_w_1_120_s_0_280 = 5.65e-12
+ mcm4m2p1_ca_w_1_120_s_0_350 = 3.67e-05  mcm4m2p1_cc_w_1_120_s_0_350 = 7.73e-11  mcm4m2p1_cf_w_1_120_s_0_350 = 6.86e-12
+ mcm4m2p1_ca_w_1_120_s_0_420 = 3.67e-05  mcm4m2p1_cc_w_1_120_s_0_420 = 6.84e-11  mcm4m2p1_cf_w_1_120_s_0_420 = 8.05e-12
+ mcm4m2p1_ca_w_1_120_s_0_560 = 3.67e-05  mcm4m2p1_cc_w_1_120_s_0_560 = 5.51e-11  mcm4m2p1_cf_w_1_120_s_0_560 = 1.04e-11
+ mcm4m2p1_ca_w_1_120_s_0_840 = 3.67e-05  mcm4m2p1_cc_w_1_120_s_0_840 = 3.92e-11  mcm4m2p1_cf_w_1_120_s_0_840 = 1.48e-11
+ mcm4m2p1_ca_w_1_120_s_1_540 = 3.67e-05  mcm4m2p1_cc_w_1_120_s_1_540 = 2.03e-11  mcm4m2p1_cf_w_1_120_s_1_540 = 2.36e-11
+ mcm4m2p1_ca_w_1_120_s_3_500 = 3.67e-05  mcm4m2p1_cc_w_1_120_s_3_500 = 4.30e-12  mcm4m2p1_cf_w_1_120_s_3_500 = 3.55e-11
+ mcm4m2l1_ca_w_0_140_s_0_140 = 4.64e-05  mcm4m2l1_cc_w_0_140_s_0_140 = 8.48e-11  mcm4m2l1_cf_w_0_140_s_0_140 = 3.88e-12
+ mcm4m2l1_ca_w_0_140_s_0_175 = 4.64e-05  mcm4m2l1_cc_w_0_140_s_0_175 = 8.39e-11  mcm4m2l1_cf_w_0_140_s_0_175 = 4.68e-12
+ mcm4m2l1_ca_w_0_140_s_0_210 = 4.64e-05  mcm4m2l1_cc_w_0_140_s_0_210 = 8.05e-11  mcm4m2l1_cf_w_0_140_s_0_210 = 5.51e-12
+ mcm4m2l1_ca_w_0_140_s_0_280 = 4.64e-05  mcm4m2l1_cc_w_0_140_s_0_280 = 7.18e-11  mcm4m2l1_cf_w_0_140_s_0_280 = 7.04e-12
+ mcm4m2l1_ca_w_0_140_s_0_350 = 4.64e-05  mcm4m2l1_cc_w_0_140_s_0_350 = 6.27e-11  mcm4m2l1_cf_w_0_140_s_0_350 = 8.55e-12
+ mcm4m2l1_ca_w_0_140_s_0_420 = 4.64e-05  mcm4m2l1_cc_w_0_140_s_0_420 = 5.44e-11  mcm4m2l1_cf_w_0_140_s_0_420 = 1.01e-11
+ mcm4m2l1_ca_w_0_140_s_0_560 = 4.64e-05  mcm4m2l1_cc_w_0_140_s_0_560 = 4.34e-11  mcm4m2l1_cf_w_0_140_s_0_560 = 1.29e-11
+ mcm4m2l1_ca_w_0_140_s_0_840 = 4.64e-05  mcm4m2l1_cc_w_0_140_s_0_840 = 2.98e-11  mcm4m2l1_cf_w_0_140_s_0_840 = 1.79e-11
+ mcm4m2l1_ca_w_0_140_s_1_540 = 4.64e-05  mcm4m2l1_cc_w_0_140_s_1_540 = 1.39e-11  mcm4m2l1_cf_w_0_140_s_1_540 = 2.73e-11
+ mcm4m2l1_ca_w_0_140_s_3_500 = 4.64e-05  mcm4m2l1_cc_w_0_140_s_3_500 = 2.19e-12  mcm4m2l1_cf_w_0_140_s_3_500 = 3.71e-11
+ mcm4m2l1_ca_w_1_120_s_0_140 = 4.64e-05  mcm4m2l1_cc_w_1_120_s_0_140 = 1.03e-10  mcm4m2l1_cf_w_1_120_s_0_140 = 3.91e-12
+ mcm4m2l1_ca_w_1_120_s_0_175 = 4.64e-05  mcm4m2l1_cc_w_1_120_s_0_175 = 1.00e-10  mcm4m2l1_cf_w_1_120_s_0_175 = 4.71e-12
+ mcm4m2l1_ca_w_1_120_s_0_210 = 4.64e-05  mcm4m2l1_cc_w_1_120_s_0_210 = 9.57e-11  mcm4m2l1_cf_w_1_120_s_0_210 = 5.50e-12
+ mcm4m2l1_ca_w_1_120_s_0_280 = 4.64e-05  mcm4m2l1_cc_w_1_120_s_0_280 = 8.46e-11  mcm4m2l1_cf_w_1_120_s_0_280 = 7.07e-12
+ mcm4m2l1_ca_w_1_120_s_0_350 = 4.64e-05  mcm4m2l1_cc_w_1_120_s_0_350 = 7.37e-11  mcm4m2l1_cf_w_1_120_s_0_350 = 8.60e-12
+ mcm4m2l1_ca_w_1_120_s_0_420 = 4.64e-05  mcm4m2l1_cc_w_1_120_s_0_420 = 6.45e-11  mcm4m2l1_cf_w_1_120_s_0_420 = 1.01e-11
+ mcm4m2l1_ca_w_1_120_s_0_560 = 4.64e-05  mcm4m2l1_cc_w_1_120_s_0_560 = 5.11e-11  mcm4m2l1_cf_w_1_120_s_0_560 = 1.30e-11
+ mcm4m2l1_ca_w_1_120_s_0_840 = 4.64e-05  mcm4m2l1_cc_w_1_120_s_0_840 = 3.51e-11  mcm4m2l1_cf_w_1_120_s_0_840 = 1.82e-11
+ mcm4m2l1_ca_w_1_120_s_1_540 = 4.64e-05  mcm4m2l1_cc_w_1_120_s_1_540 = 1.66e-11  mcm4m2l1_cf_w_1_120_s_1_540 = 2.82e-11
+ mcm4m2l1_ca_w_1_120_s_3_500 = 4.64e-05  mcm4m2l1_cc_w_1_120_s_3_500 = 2.73e-12  mcm4m2l1_cf_w_1_120_s_3_500 = 3.96e-11
+ mcm4m2m1_ca_w_0_140_s_0_140 = 9.81e-05  mcm4m2m1_cc_w_0_140_s_0_140 = 7.97e-11  mcm4m2m1_cf_w_0_140_s_0_140 = 7.93e-12
+ mcm4m2m1_ca_w_0_140_s_0_175 = 9.81e-05  mcm4m2m1_cc_w_0_140_s_0_175 = 7.81e-11  mcm4m2m1_cf_w_0_140_s_0_175 = 9.63e-12
+ mcm4m2m1_ca_w_0_140_s_0_210 = 9.81e-05  mcm4m2m1_cc_w_0_140_s_0_210 = 7.44e-11  mcm4m2m1_cf_w_0_140_s_0_210 = 1.13e-11
+ mcm4m2m1_ca_w_0_140_s_0_280 = 9.81e-05  mcm4m2m1_cc_w_0_140_s_0_280 = 6.45e-11  mcm4m2m1_cf_w_0_140_s_0_280 = 1.44e-11
+ mcm4m2m1_ca_w_0_140_s_0_350 = 9.81e-05  mcm4m2m1_cc_w_0_140_s_0_350 = 5.51e-11  mcm4m2m1_cf_w_0_140_s_0_350 = 1.74e-11
+ mcm4m2m1_ca_w_0_140_s_0_420 = 9.81e-05  mcm4m2m1_cc_w_0_140_s_0_420 = 4.65e-11  mcm4m2m1_cf_w_0_140_s_0_420 = 2.01e-11
+ mcm4m2m1_ca_w_0_140_s_0_560 = 9.81e-05  mcm4m2m1_cc_w_0_140_s_0_560 = 3.49e-11  mcm4m2m1_cf_w_0_140_s_0_560 = 2.53e-11
+ mcm4m2m1_ca_w_0_140_s_0_840 = 9.81e-05  mcm4m2m1_cc_w_0_140_s_0_840 = 2.13e-11  mcm4m2m1_cf_w_0_140_s_0_840 = 3.32e-11
+ mcm4m2m1_ca_w_0_140_s_1_540 = 9.81e-05  mcm4m2m1_cc_w_0_140_s_1_540 = 7.44e-12  mcm4m2m1_cf_w_0_140_s_1_540 = 4.41e-11
+ mcm4m2m1_ca_w_0_140_s_3_500 = 9.81e-05  mcm4m2m1_cc_w_0_140_s_3_500 = 6.75e-13  mcm4m2m1_cf_w_0_140_s_3_500 = 5.08e-11
+ mcm4m2m1_ca_w_1_120_s_0_140 = 9.81e-05  mcm4m2m1_cc_w_1_120_s_0_140 = 9.20e-11  mcm4m2m1_cf_w_1_120_s_0_140 = 7.94e-12
+ mcm4m2m1_ca_w_1_120_s_0_175 = 9.81e-05  mcm4m2m1_cc_w_1_120_s_0_175 = 8.95e-11  mcm4m2m1_cf_w_1_120_s_0_175 = 9.64e-12
+ mcm4m2m1_ca_w_1_120_s_0_210 = 9.81e-05  mcm4m2m1_cc_w_1_120_s_0_210 = 8.48e-11  mcm4m2m1_cf_w_1_120_s_0_210 = 1.13e-11
+ mcm4m2m1_ca_w_1_120_s_0_280 = 9.81e-05  mcm4m2m1_cc_w_1_120_s_0_280 = 7.36e-11  mcm4m2m1_cf_w_1_120_s_0_280 = 1.44e-11
+ mcm4m2m1_ca_w_1_120_s_0_350 = 9.81e-05  mcm4m2m1_cc_w_1_120_s_0_350 = 6.26e-11  mcm4m2m1_cf_w_1_120_s_0_350 = 1.74e-11
+ mcm4m2m1_ca_w_1_120_s_0_420 = 9.81e-05  mcm4m2m1_cc_w_1_120_s_0_420 = 5.35e-11  mcm4m2m1_cf_w_1_120_s_0_420 = 2.03e-11
+ mcm4m2m1_ca_w_1_120_s_0_560 = 9.81e-05  mcm4m2m1_cc_w_1_120_s_0_560 = 4.05e-11  mcm4m2m1_cf_w_1_120_s_0_560 = 2.53e-11
+ mcm4m2m1_ca_w_1_120_s_0_840 = 9.81e-05  mcm4m2m1_cc_w_1_120_s_0_840 = 2.51e-11  mcm4m2m1_cf_w_1_120_s_0_840 = 3.36e-11
+ mcm4m2m1_ca_w_1_120_s_1_540 = 9.81e-05  mcm4m2m1_cc_w_1_120_s_1_540 = 9.42e-12  mcm4m2m1_cf_w_1_120_s_1_540 = 4.55e-11
+ mcm4m2m1_ca_w_1_120_s_3_500 = 9.81e-05  mcm4m2m1_cc_w_1_120_s_3_500 = 9.00e-13  mcm4m2m1_cf_w_1_120_s_3_500 = 5.36e-11
+ mcm5m2f_ca_w_0_140_s_0_140 = 2.41e-05  mcm5m2f_cc_w_0_140_s_0_140 = 8.80e-11  mcm5m2f_cf_w_0_140_s_0_140 = 2.04e-12
+ mcm5m2f_ca_w_0_140_s_0_175 = 2.41e-05  mcm5m2f_cc_w_0_140_s_0_175 = 8.61e-11  mcm5m2f_cf_w_0_140_s_0_175 = 2.45e-12
+ mcm5m2f_ca_w_0_140_s_0_210 = 2.41e-05  mcm5m2f_cc_w_0_140_s_0_210 = 8.34e-11  mcm5m2f_cf_w_0_140_s_0_210 = 2.90e-12
+ mcm5m2f_ca_w_0_140_s_0_280 = 2.41e-05  mcm5m2f_cc_w_0_140_s_0_280 = 7.56e-11  mcm5m2f_cf_w_0_140_s_0_280 = 3.70e-12
+ mcm5m2f_ca_w_0_140_s_0_350 = 2.41e-05  mcm5m2f_cc_w_0_140_s_0_350 = 6.70e-11  mcm5m2f_cf_w_0_140_s_0_350 = 4.51e-12
+ mcm5m2f_ca_w_0_140_s_0_420 = 2.41e-05  mcm5m2f_cc_w_0_140_s_0_420 = 5.91e-11  mcm5m2f_cf_w_0_140_s_0_420 = 5.35e-12
+ mcm5m2f_ca_w_0_140_s_0_560 = 2.41e-05  mcm5m2f_cc_w_0_140_s_0_560 = 4.91e-11  mcm5m2f_cf_w_0_140_s_0_560 = 6.93e-12
+ mcm5m2f_ca_w_0_140_s_0_840 = 2.41e-05  mcm5m2f_cc_w_0_140_s_0_840 = 3.68e-11  mcm5m2f_cf_w_0_140_s_0_840 = 9.85e-12
+ mcm5m2f_ca_w_0_140_s_1_540 = 2.41e-05  mcm5m2f_cc_w_0_140_s_1_540 = 2.17e-11  mcm5m2f_cf_w_0_140_s_1_540 = 1.61e-11
+ mcm5m2f_ca_w_0_140_s_3_500 = 2.41e-05  mcm5m2f_cc_w_0_140_s_3_500 = 6.93e-12  mcm5m2f_cf_w_0_140_s_3_500 = 2.62e-11
+ mcm5m2f_ca_w_1_120_s_0_140 = 2.41e-05  mcm5m2f_cc_w_1_120_s_0_140 = 1.12e-10  mcm5m2f_cf_w_1_120_s_0_140 = 2.06e-12
+ mcm5m2f_ca_w_1_120_s_0_175 = 2.41e-05  mcm5m2f_cc_w_1_120_s_0_175 = 1.10e-10  mcm5m2f_cf_w_1_120_s_0_175 = 2.47e-12
+ mcm5m2f_ca_w_1_120_s_0_210 = 2.41e-05  mcm5m2f_cc_w_1_120_s_0_210 = 1.06e-10  mcm5m2f_cf_w_1_120_s_0_210 = 2.89e-12
+ mcm5m2f_ca_w_1_120_s_0_280 = 2.41e-05  mcm5m2f_cc_w_1_120_s_0_280 = 9.37e-11  mcm5m2f_cf_w_1_120_s_0_280 = 3.72e-12
+ mcm5m2f_ca_w_1_120_s_0_350 = 2.41e-05  mcm5m2f_cc_w_1_120_s_0_350 = 8.37e-11  mcm5m2f_cf_w_1_120_s_0_350 = 4.54e-12
+ mcm5m2f_ca_w_1_120_s_0_420 = 2.41e-05  mcm5m2f_cc_w_1_120_s_0_420 = 7.48e-11  mcm5m2f_cf_w_1_120_s_0_420 = 5.35e-12
+ mcm5m2f_ca_w_1_120_s_0_560 = 2.41e-05  mcm5m2f_cc_w_1_120_s_0_560 = 6.20e-11  mcm5m2f_cf_w_1_120_s_0_560 = 6.93e-12
+ mcm5m2f_ca_w_1_120_s_0_840 = 2.41e-05  mcm5m2f_cc_w_1_120_s_0_840 = 4.63e-11  mcm5m2f_cf_w_1_120_s_0_840 = 9.96e-12
+ mcm5m2f_ca_w_1_120_s_1_540 = 2.41e-05  mcm5m2f_cc_w_1_120_s_1_540 = 2.76e-11  mcm5m2f_cf_w_1_120_s_1_540 = 1.66e-11
+ mcm5m2f_ca_w_1_120_s_3_500 = 2.41e-05  mcm5m2f_cc_w_1_120_s_3_500 = 9.07e-12  mcm5m2f_cf_w_1_120_s_3_500 = 2.82e-11
+ mcm5m2d_ca_w_0_140_s_0_140 = 2.69e-05  mcm5m2d_cc_w_0_140_s_0_140 = 8.78e-11  mcm5m2d_cf_w_0_140_s_0_140 = 2.28e-12
+ mcm5m2d_ca_w_0_140_s_0_175 = 2.69e-05  mcm5m2d_cc_w_0_140_s_0_175 = 8.59e-11  mcm5m2d_cf_w_0_140_s_0_175 = 2.74e-12
+ mcm5m2d_ca_w_0_140_s_0_210 = 2.69e-05  mcm5m2d_cc_w_0_140_s_0_210 = 8.28e-11  mcm5m2d_cf_w_0_140_s_0_210 = 3.23e-12
+ mcm5m2d_ca_w_0_140_s_0_280 = 2.69e-05  mcm5m2d_cc_w_0_140_s_0_280 = 7.52e-11  mcm5m2d_cf_w_0_140_s_0_280 = 4.13e-12
+ mcm5m2d_ca_w_0_140_s_0_350 = 2.69e-05  mcm5m2d_cc_w_0_140_s_0_350 = 6.64e-11  mcm5m2d_cf_w_0_140_s_0_350 = 5.04e-12
+ mcm5m2d_ca_w_0_140_s_0_420 = 2.69e-05  mcm5m2d_cc_w_0_140_s_0_420 = 5.86e-11  mcm5m2d_cf_w_0_140_s_0_420 = 5.96e-12
+ mcm5m2d_ca_w_0_140_s_0_560 = 2.69e-05  mcm5m2d_cc_w_0_140_s_0_560 = 4.83e-11  mcm5m2d_cf_w_0_140_s_0_560 = 7.71e-12
+ mcm5m2d_ca_w_0_140_s_0_840 = 2.69e-05  mcm5m2d_cc_w_0_140_s_0_840 = 3.58e-11  mcm5m2d_cf_w_0_140_s_0_840 = 1.09e-11
+ mcm5m2d_ca_w_0_140_s_1_540 = 2.69e-05  mcm5m2d_cc_w_0_140_s_1_540 = 2.05e-11  mcm5m2d_cf_w_0_140_s_1_540 = 1.77e-11
+ mcm5m2d_ca_w_0_140_s_3_500 = 2.69e-05  mcm5m2d_cc_w_0_140_s_3_500 = 6.03e-12  mcm5m2d_cf_w_0_140_s_3_500 = 2.80e-11
+ mcm5m2d_ca_w_1_120_s_0_140 = 2.69e-05  mcm5m2d_cc_w_1_120_s_0_140 = 1.11e-10  mcm5m2d_cf_w_1_120_s_0_140 = 2.30e-12
+ mcm5m2d_ca_w_1_120_s_0_175 = 2.69e-05  mcm5m2d_cc_w_1_120_s_0_175 = 1.09e-10  mcm5m2d_cf_w_1_120_s_0_175 = 2.77e-12
+ mcm5m2d_ca_w_1_120_s_0_210 = 2.69e-05  mcm5m2d_cc_w_1_120_s_0_210 = 1.04e-10  mcm5m2d_cf_w_1_120_s_0_210 = 3.23e-12
+ mcm5m2d_ca_w_1_120_s_0_280 = 2.69e-05  mcm5m2d_cc_w_1_120_s_0_280 = 9.23e-11  mcm5m2d_cf_w_1_120_s_0_280 = 4.15e-12
+ mcm5m2d_ca_w_1_120_s_0_350 = 2.69e-05  mcm5m2d_cc_w_1_120_s_0_350 = 8.23e-11  mcm5m2d_cf_w_1_120_s_0_350 = 5.07e-12
+ mcm5m2d_ca_w_1_120_s_0_420 = 2.69e-05  mcm5m2d_cc_w_1_120_s_0_420 = 7.33e-11  mcm5m2d_cf_w_1_120_s_0_420 = 5.97e-12
+ mcm5m2d_ca_w_1_120_s_0_560 = 2.69e-05  mcm5m2d_cc_w_1_120_s_0_560 = 6.05e-11  mcm5m2d_cf_w_1_120_s_0_560 = 7.73e-12
+ mcm5m2d_ca_w_1_120_s_0_840 = 2.69e-05  mcm5m2d_cc_w_1_120_s_0_840 = 4.46e-11  mcm5m2d_cf_w_1_120_s_0_840 = 1.11e-11
+ mcm5m2d_ca_w_1_120_s_1_540 = 2.69e-05  mcm5m2d_cc_w_1_120_s_1_540 = 2.59e-11  mcm5m2d_cf_w_1_120_s_1_540 = 1.82e-11
+ mcm5m2d_ca_w_1_120_s_3_500 = 2.69e-05  mcm5m2d_cc_w_1_120_s_3_500 = 7.88e-12  mcm5m2d_cf_w_1_120_s_3_500 = 3.01e-11
+ mcm5m2p1_ca_w_0_140_s_0_140 = 2.90e-05  mcm5m2p1_cc_w_0_140_s_0_140 = 8.76e-11  mcm5m2p1_cf_w_0_140_s_0_140 = 2.46e-12
+ mcm5m2p1_ca_w_0_140_s_0_175 = 2.90e-05  mcm5m2p1_cc_w_0_140_s_0_175 = 8.55e-11  mcm5m2p1_cf_w_0_140_s_0_175 = 2.95e-12
+ mcm5m2p1_ca_w_0_140_s_0_210 = 2.90e-05  mcm5m2p1_cc_w_0_140_s_0_210 = 8.25e-11  mcm5m2p1_cf_w_0_140_s_0_210 = 3.49e-12
+ mcm5m2p1_ca_w_0_140_s_0_280 = 2.90e-05  mcm5m2p1_cc_w_0_140_s_0_280 = 7.48e-11  mcm5m2p1_cf_w_0_140_s_0_280 = 4.46e-12
+ mcm5m2p1_ca_w_0_140_s_0_350 = 2.90e-05  mcm5m2p1_cc_w_0_140_s_0_350 = 6.60e-11  mcm5m2p1_cf_w_0_140_s_0_350 = 5.43e-12
+ mcm5m2p1_ca_w_0_140_s_0_420 = 2.90e-05  mcm5m2p1_cc_w_0_140_s_0_420 = 5.81e-11  mcm5m2p1_cf_w_0_140_s_0_420 = 6.43e-12
+ mcm5m2p1_ca_w_0_140_s_0_560 = 2.90e-05  mcm5m2p1_cc_w_0_140_s_0_560 = 4.77e-11  mcm5m2p1_cf_w_0_140_s_0_560 = 8.30e-12
+ mcm5m2p1_ca_w_0_140_s_0_840 = 2.90e-05  mcm5m2p1_cc_w_0_140_s_0_840 = 3.50e-11  mcm5m2p1_cf_w_0_140_s_0_840 = 1.17e-11
+ mcm5m2p1_ca_w_0_140_s_1_540 = 2.90e-05  mcm5m2p1_cc_w_0_140_s_1_540 = 1.97e-11  mcm5m2p1_cf_w_0_140_s_1_540 = 1.88e-11
+ mcm5m2p1_ca_w_0_140_s_3_500 = 2.90e-05  mcm5m2p1_cc_w_0_140_s_3_500 = 5.47e-12  mcm5m2p1_cf_w_0_140_s_3_500 = 2.92e-11
+ mcm5m2p1_ca_w_1_120_s_0_140 = 2.90e-05  mcm5m2p1_cc_w_1_120_s_0_140 = 1.10e-10  mcm5m2p1_cf_w_1_120_s_0_140 = 2.50e-12
+ mcm5m2p1_ca_w_1_120_s_0_175 = 2.90e-05  mcm5m2p1_cc_w_1_120_s_0_175 = 1.08e-10  mcm5m2p1_cf_w_1_120_s_0_175 = 3.00e-12
+ mcm5m2p1_ca_w_1_120_s_0_210 = 2.90e-05  mcm5m2p1_cc_w_1_120_s_0_210 = 1.03e-10  mcm5m2p1_cf_w_1_120_s_0_210 = 3.50e-12
+ mcm5m2p1_ca_w_1_120_s_0_280 = 2.90e-05  mcm5m2p1_cc_w_1_120_s_0_280 = 9.13e-11  mcm5m2p1_cf_w_1_120_s_0_280 = 4.50e-12
+ mcm5m2p1_ca_w_1_120_s_0_350 = 2.90e-05  mcm5m2p1_cc_w_1_120_s_0_350 = 8.12e-11  mcm5m2p1_cf_w_1_120_s_0_350 = 5.48e-12
+ mcm5m2p1_ca_w_1_120_s_0_420 = 2.90e-05  mcm5m2p1_cc_w_1_120_s_0_420 = 7.25e-11  mcm5m2p1_cf_w_1_120_s_0_420 = 6.45e-12
+ mcm5m2p1_ca_w_1_120_s_0_560 = 2.90e-05  mcm5m2p1_cc_w_1_120_s_0_560 = 5.94e-11  mcm5m2p1_cf_w_1_120_s_0_560 = 8.33e-12
+ mcm5m2p1_ca_w_1_120_s_0_840 = 2.90e-05  mcm5m2p1_cc_w_1_120_s_0_840 = 4.36e-11  mcm5m2p1_cf_w_1_120_s_0_840 = 1.19e-11
+ mcm5m2p1_ca_w_1_120_s_1_540 = 2.90e-05  mcm5m2p1_cc_w_1_120_s_1_540 = 2.47e-11  mcm5m2p1_cf_w_1_120_s_1_540 = 1.95e-11
+ mcm5m2p1_ca_w_1_120_s_3_500 = 2.90e-05  mcm5m2p1_cc_w_1_120_s_3_500 = 7.16e-12  mcm5m2p1_cf_w_1_120_s_3_500 = 3.15e-11
+ mcm5m2l1_ca_w_0_140_s_0_140 = 3.87e-05  mcm5m2l1_cc_w_0_140_s_0_140 = 8.58e-11  mcm5m2l1_cf_w_0_140_s_0_140 = 3.25e-12
+ mcm5m2l1_ca_w_0_140_s_0_175 = 3.87e-05  mcm5m2l1_cc_w_0_140_s_0_175 = 8.47e-11  mcm5m2l1_cf_w_0_140_s_0_175 = 3.92e-12
+ mcm5m2l1_ca_w_0_140_s_0_210 = 3.87e-05  mcm5m2l1_cc_w_0_140_s_0_210 = 8.11e-11  mcm5m2l1_cf_w_0_140_s_0_210 = 4.61e-12
+ mcm5m2l1_ca_w_0_140_s_0_280 = 3.87e-05  mcm5m2l1_cc_w_0_140_s_0_280 = 7.32e-11  mcm5m2l1_cf_w_0_140_s_0_280 = 5.90e-12
+ mcm5m2l1_ca_w_0_140_s_0_350 = 3.87e-05  mcm5m2l1_cc_w_0_140_s_0_350 = 6.43e-11  mcm5m2l1_cf_w_0_140_s_0_350 = 7.18e-12
+ mcm5m2l1_ca_w_0_140_s_0_420 = 3.87e-05  mcm5m2l1_cc_w_0_140_s_0_420 = 5.62e-11  mcm5m2l1_cf_w_0_140_s_0_420 = 8.48e-12
+ mcm5m2l1_ca_w_0_140_s_0_560 = 3.87e-05  mcm5m2l1_cc_w_0_140_s_0_560 = 4.53e-11  mcm5m2l1_cf_w_0_140_s_0_560 = 1.09e-11
+ mcm5m2l1_ca_w_0_140_s_0_840 = 3.87e-05  mcm5m2l1_cc_w_0_140_s_0_840 = 3.22e-11  mcm5m2l1_cf_w_0_140_s_0_840 = 1.52e-11
+ mcm5m2l1_ca_w_0_140_s_1_540 = 3.87e-05  mcm5m2l1_cc_w_0_140_s_1_540 = 1.67e-11  mcm5m2l1_cf_w_0_140_s_1_540 = 2.37e-11
+ mcm5m2l1_ca_w_0_140_s_3_500 = 3.87e-05  mcm5m2l1_cc_w_0_140_s_3_500 = 3.76e-12  mcm5m2l1_cf_w_0_140_s_3_500 = 3.40e-11
+ mcm5m2l1_ca_w_1_120_s_0_140 = 3.87e-05  mcm5m2l1_cc_w_1_120_s_0_140 = 1.06e-10  mcm5m2l1_cf_w_1_120_s_0_140 = 3.28e-12
+ mcm5m2l1_ca_w_1_120_s_0_175 = 3.87e-05  mcm5m2l1_cc_w_1_120_s_0_175 = 1.04e-10  mcm5m2l1_cf_w_1_120_s_0_175 = 3.95e-12
+ mcm5m2l1_ca_w_1_120_s_0_210 = 3.87e-05  mcm5m2l1_cc_w_1_120_s_0_210 = 9.93e-11  mcm5m2l1_cf_w_1_120_s_0_210 = 4.61e-12
+ mcm5m2l1_ca_w_1_120_s_0_280 = 3.87e-05  mcm5m2l1_cc_w_1_120_s_0_280 = 8.81e-11  mcm5m2l1_cf_w_1_120_s_0_280 = 5.95e-12
+ mcm5m2l1_ca_w_1_120_s_0_350 = 3.87e-05  mcm5m2l1_cc_w_1_120_s_0_350 = 7.73e-11  mcm5m2l1_cf_w_1_120_s_0_350 = 7.22e-12
+ mcm5m2l1_ca_w_1_120_s_0_420 = 3.87e-05  mcm5m2l1_cc_w_1_120_s_0_420 = 6.85e-11  mcm5m2l1_cf_w_1_120_s_0_420 = 8.48e-12
+ mcm5m2l1_ca_w_1_120_s_0_560 = 3.87e-05  mcm5m2l1_cc_w_1_120_s_0_560 = 5.53e-11  mcm5m2l1_cf_w_1_120_s_0_560 = 1.09e-11
+ mcm5m2l1_ca_w_1_120_s_0_840 = 3.87e-05  mcm5m2l1_cc_w_1_120_s_0_840 = 3.95e-11  mcm5m2l1_cf_w_1_120_s_0_840 = 1.54e-11
+ mcm5m2l1_ca_w_1_120_s_1_540 = 3.87e-05  mcm5m2l1_cc_w_1_120_s_1_540 = 2.09e-11  mcm5m2l1_cf_w_1_120_s_1_540 = 2.44e-11
+ mcm5m2l1_ca_w_1_120_s_3_500 = 3.87e-05  mcm5m2l1_cc_w_1_120_s_3_500 = 5.07e-12  mcm5m2l1_cf_w_1_120_s_3_500 = 3.65e-11
+ mcm5m2m1_ca_w_0_140_s_0_140 = 9.05e-05  mcm5m2m1_cc_w_0_140_s_0_140 = 8.07e-11  mcm5m2m1_cf_w_0_140_s_0_140 = 7.30e-12
+ mcm5m2m1_ca_w_0_140_s_0_175 = 9.05e-05  mcm5m2m1_cc_w_0_140_s_0_175 = 7.91e-11  mcm5m2m1_cf_w_0_140_s_0_175 = 8.87e-12
+ mcm5m2m1_ca_w_0_140_s_0_210 = 9.05e-05  mcm5m2m1_cc_w_0_140_s_0_210 = 7.51e-11  mcm5m2m1_cf_w_0_140_s_0_210 = 1.04e-11
+ mcm5m2m1_ca_w_0_140_s_0_280 = 9.05e-05  mcm5m2m1_cc_w_0_140_s_0_280 = 6.62e-11  mcm5m2m1_cf_w_0_140_s_0_280 = 1.33e-11
+ mcm5m2m1_ca_w_0_140_s_0_350 = 9.05e-05  mcm5m2m1_cc_w_0_140_s_0_350 = 5.60e-11  mcm5m2m1_cf_w_0_140_s_0_350 = 1.60e-11
+ mcm5m2m1_ca_w_0_140_s_0_420 = 9.05e-05  mcm5m2m1_cc_w_0_140_s_0_420 = 4.83e-11  mcm5m2m1_cf_w_0_140_s_0_420 = 1.86e-11
+ mcm5m2m1_ca_w_0_140_s_0_560 = 9.05e-05  mcm5m2m1_cc_w_0_140_s_0_560 = 3.68e-11  mcm5m2m1_cf_w_0_140_s_0_560 = 2.33e-11
+ mcm5m2m1_ca_w_0_140_s_0_840 = 9.05e-05  mcm5m2m1_cc_w_0_140_s_0_840 = 2.35e-11  mcm5m2m1_cf_w_0_140_s_0_840 = 3.08e-11
+ mcm5m2m1_ca_w_0_140_s_1_540 = 9.05e-05  mcm5m2m1_cc_w_0_140_s_1_540 = 9.52e-12  mcm5m2m1_cf_w_0_140_s_1_540 = 4.16e-11
+ mcm5m2m1_ca_w_0_140_s_3_500 = 9.05e-05  mcm5m2m1_cc_w_0_140_s_3_500 = 1.43e-12  mcm5m2m1_cf_w_0_140_s_3_500 = 4.92e-11
+ mcm5m2m1_ca_w_1_120_s_0_140 = 9.05e-05  mcm5m2m1_cc_w_1_120_s_0_140 = 9.56e-11  mcm5m2m1_cf_w_1_120_s_0_140 = 7.30e-12
+ mcm5m2m1_ca_w_1_120_s_0_175 = 9.05e-05  mcm5m2m1_cc_w_1_120_s_0_175 = 9.31e-11  mcm5m2m1_cf_w_1_120_s_0_175 = 8.88e-12
+ mcm5m2m1_ca_w_1_120_s_0_210 = 9.05e-05  mcm5m2m1_cc_w_1_120_s_0_210 = 8.84e-11  mcm5m2m1_cf_w_1_120_s_0_210 = 1.04e-11
+ mcm5m2m1_ca_w_1_120_s_0_280 = 9.05e-05  mcm5m2m1_cc_w_1_120_s_0_280 = 7.73e-11  mcm5m2m1_cf_w_1_120_s_0_280 = 1.33e-11
+ mcm5m2m1_ca_w_1_120_s_0_350 = 9.05e-05  mcm5m2m1_cc_w_1_120_s_0_350 = 6.64e-11  mcm5m2m1_cf_w_1_120_s_0_350 = 1.60e-11
+ mcm5m2m1_ca_w_1_120_s_0_420 = 9.05e-05  mcm5m2m1_cc_w_1_120_s_0_420 = 5.76e-11  mcm5m2m1_cf_w_1_120_s_0_420 = 1.87e-11
+ mcm5m2m1_ca_w_1_120_s_0_560 = 9.05e-05  mcm5m2m1_cc_w_1_120_s_0_560 = 4.46e-11  mcm5m2m1_cf_w_1_120_s_0_560 = 2.34e-11
+ mcm5m2m1_ca_w_1_120_s_0_840 = 9.05e-05  mcm5m2m1_cc_w_1_120_s_0_840 = 2.94e-11  mcm5m2m1_cf_w_1_120_s_0_840 = 3.10e-11
+ mcm5m2m1_ca_w_1_120_s_1_540 = 9.05e-05  mcm5m2m1_cc_w_1_120_s_1_540 = 1.30e-11  mcm5m2m1_cf_w_1_120_s_1_540 = 4.28e-11
+ mcm5m2m1_ca_w_1_120_s_3_500 = 9.05e-05  mcm5m2m1_cc_w_1_120_s_3_500 = 2.25e-12  mcm5m2m1_cf_w_1_120_s_3_500 = 5.27e-11
+ mcrdlm2f_ca_w_0_140_s_0_140 = 1.66e-05  mcrdlm2f_cc_w_0_140_s_0_140 = 8.85e-11  mcrdlm2f_cf_w_0_140_s_0_140 = 1.41e-12
+ mcrdlm2f_ca_w_0_140_s_0_175 = 1.66e-05  mcrdlm2f_cc_w_0_140_s_0_175 = 8.70e-11  mcrdlm2f_cf_w_0_140_s_0_175 = 1.70e-12
+ mcrdlm2f_ca_w_0_140_s_0_210 = 1.66e-05  mcrdlm2f_cc_w_0_140_s_0_210 = 8.42e-11  mcrdlm2f_cf_w_0_140_s_0_210 = 2.00e-12
+ mcrdlm2f_ca_w_0_140_s_0_280 = 1.66e-05  mcrdlm2f_cc_w_0_140_s_0_280 = 7.68e-11  mcrdlm2f_cf_w_0_140_s_0_280 = 2.57e-12
+ mcrdlm2f_ca_w_0_140_s_0_350 = 1.66e-05  mcrdlm2f_cc_w_0_140_s_0_350 = 6.81e-11  mcrdlm2f_cf_w_0_140_s_0_350 = 3.12e-12
+ mcrdlm2f_ca_w_0_140_s_0_420 = 1.66e-05  mcrdlm2f_cc_w_0_140_s_0_420 = 6.09e-11  mcrdlm2f_cf_w_0_140_s_0_420 = 3.71e-12
+ mcrdlm2f_ca_w_0_140_s_0_560 = 1.66e-05  mcrdlm2f_cc_w_0_140_s_0_560 = 5.11e-11  mcrdlm2f_cf_w_0_140_s_0_560 = 4.80e-12
+ mcrdlm2f_ca_w_0_140_s_0_840 = 1.66e-05  mcrdlm2f_cc_w_0_140_s_0_840 = 3.96e-11  mcrdlm2f_cf_w_0_140_s_0_840 = 6.88e-12
+ mcrdlm2f_ca_w_0_140_s_1_540 = 1.66e-05  mcrdlm2f_cc_w_0_140_s_1_540 = 2.57e-11  mcrdlm2f_cf_w_0_140_s_1_540 = 1.16e-11
+ mcrdlm2f_ca_w_0_140_s_3_500 = 1.66e-05  mcrdlm2f_cc_w_0_140_s_3_500 = 1.14e-11  mcrdlm2f_cf_w_0_140_s_3_500 = 2.03e-11
+ mcrdlm2f_ca_w_1_120_s_0_140 = 1.66e-05  mcrdlm2f_cc_w_1_120_s_0_140 = 1.17e-10  mcrdlm2f_cf_w_1_120_s_0_140 = 1.43e-12
+ mcrdlm2f_ca_w_1_120_s_0_175 = 1.66e-05  mcrdlm2f_cc_w_1_120_s_0_175 = 1.14e-10  mcrdlm2f_cf_w_1_120_s_0_175 = 1.72e-12
+ mcrdlm2f_ca_w_1_120_s_0_210 = 1.66e-05  mcrdlm2f_cc_w_1_120_s_0_210 = 1.09e-10  mcrdlm2f_cf_w_1_120_s_0_210 = 2.01e-12
+ mcrdlm2f_ca_w_1_120_s_0_280 = 1.66e-05  mcrdlm2f_cc_w_1_120_s_0_280 = 9.81e-11  mcrdlm2f_cf_w_1_120_s_0_280 = 2.58e-12
+ mcrdlm2f_ca_w_1_120_s_0_350 = 1.66e-05  mcrdlm2f_cc_w_1_120_s_0_350 = 8.84e-11  mcrdlm2f_cf_w_1_120_s_0_350 = 3.15e-12
+ mcrdlm2f_ca_w_1_120_s_0_420 = 1.66e-05  mcrdlm2f_cc_w_1_120_s_0_420 = 7.93e-11  mcrdlm2f_cf_w_1_120_s_0_420 = 3.71e-12
+ mcrdlm2f_ca_w_1_120_s_0_560 = 1.66e-05  mcrdlm2f_cc_w_1_120_s_0_560 = 6.68e-11  mcrdlm2f_cf_w_1_120_s_0_560 = 4.81e-12
+ mcrdlm2f_ca_w_1_120_s_0_840 = 1.66e-05  mcrdlm2f_cc_w_1_120_s_0_840 = 5.20e-11  mcrdlm2f_cf_w_1_120_s_0_840 = 6.96e-12
+ mcrdlm2f_ca_w_1_120_s_1_540 = 1.66e-05  mcrdlm2f_cc_w_1_120_s_1_540 = 3.42e-11  mcrdlm2f_cf_w_1_120_s_1_540 = 1.18e-11
+ mcrdlm2f_ca_w_1_120_s_3_500 = 1.66e-05  mcrdlm2f_cc_w_1_120_s_3_500 = 1.58e-11  mcrdlm2f_cf_w_1_120_s_3_500 = 2.17e-11
+ mcrdlm2d_ca_w_0_140_s_0_140 = 1.94e-05  mcrdlm2d_cc_w_0_140_s_0_140 = 8.81e-11  mcrdlm2d_cf_w_0_140_s_0_140 = 1.65e-12
+ mcrdlm2d_ca_w_0_140_s_0_175 = 1.94e-05  mcrdlm2d_cc_w_0_140_s_0_175 = 8.67e-11  mcrdlm2d_cf_w_0_140_s_0_175 = 1.98e-12
+ mcrdlm2d_ca_w_0_140_s_0_210 = 1.94e-05  mcrdlm2d_cc_w_0_140_s_0_210 = 8.38e-11  mcrdlm2d_cf_w_0_140_s_0_210 = 2.33e-12
+ mcrdlm2d_ca_w_0_140_s_0_280 = 1.94e-05  mcrdlm2d_cc_w_0_140_s_0_280 = 7.66e-11  mcrdlm2d_cf_w_0_140_s_0_280 = 2.99e-12
+ mcrdlm2d_ca_w_0_140_s_0_350 = 1.94e-05  mcrdlm2d_cc_w_0_140_s_0_350 = 6.75e-11  mcrdlm2d_cf_w_0_140_s_0_350 = 3.65e-12
+ mcrdlm2d_ca_w_0_140_s_0_420 = 1.94e-05  mcrdlm2d_cc_w_0_140_s_0_420 = 6.03e-11  mcrdlm2d_cf_w_0_140_s_0_420 = 4.33e-12
+ mcrdlm2d_ca_w_0_140_s_0_560 = 1.94e-05  mcrdlm2d_cc_w_0_140_s_0_560 = 5.04e-11  mcrdlm2d_cf_w_0_140_s_0_560 = 5.59e-12
+ mcrdlm2d_ca_w_0_140_s_0_840 = 1.94e-05  mcrdlm2d_cc_w_0_140_s_0_840 = 3.86e-11  mcrdlm2d_cf_w_0_140_s_0_840 = 7.98e-12
+ mcrdlm2d_ca_w_0_140_s_1_540 = 1.94e-05  mcrdlm2d_cc_w_0_140_s_1_540 = 2.44e-11  mcrdlm2d_cf_w_0_140_s_1_540 = 1.33e-11
+ mcrdlm2d_ca_w_0_140_s_3_500 = 1.94e-05  mcrdlm2d_cc_w_0_140_s_3_500 = 1.01e-11  mcrdlm2d_cf_w_0_140_s_3_500 = 2.26e-11
+ mcrdlm2d_ca_w_1_120_s_0_140 = 1.94e-05  mcrdlm2d_cc_w_1_120_s_0_140 = 1.16e-10  mcrdlm2d_cf_w_1_120_s_0_140 = 1.67e-12
+ mcrdlm2d_ca_w_1_120_s_0_175 = 1.94e-05  mcrdlm2d_cc_w_1_120_s_0_175 = 1.13e-10  mcrdlm2d_cf_w_1_120_s_0_175 = 2.02e-12
+ mcrdlm2d_ca_w_1_120_s_0_210 = 1.94e-05  mcrdlm2d_cc_w_1_120_s_0_210 = 1.08e-10  mcrdlm2d_cf_w_1_120_s_0_210 = 2.35e-12
+ mcrdlm2d_ca_w_1_120_s_0_280 = 1.94e-05  mcrdlm2d_cc_w_1_120_s_0_280 = 9.68e-11  mcrdlm2d_cf_w_1_120_s_0_280 = 3.02e-12
+ mcrdlm2d_ca_w_1_120_s_0_350 = 1.94e-05  mcrdlm2d_cc_w_1_120_s_0_350 = 8.69e-11  mcrdlm2d_cf_w_1_120_s_0_350 = 3.68e-12
+ mcrdlm2d_ca_w_1_120_s_0_420 = 1.94e-05  mcrdlm2d_cc_w_1_120_s_0_420 = 7.79e-11  mcrdlm2d_cf_w_1_120_s_0_420 = 4.34e-12
+ mcrdlm2d_ca_w_1_120_s_0_560 = 1.94e-05  mcrdlm2d_cc_w_1_120_s_0_560 = 6.54e-11  mcrdlm2d_cf_w_1_120_s_0_560 = 5.62e-12
+ mcrdlm2d_ca_w_1_120_s_0_840 = 1.94e-05  mcrdlm2d_cc_w_1_120_s_0_840 = 5.03e-11  mcrdlm2d_cf_w_1_120_s_0_840 = 8.08e-12
+ mcrdlm2d_ca_w_1_120_s_1_540 = 1.94e-05  mcrdlm2d_cc_w_1_120_s_1_540 = 3.24e-11  mcrdlm2d_cf_w_1_120_s_1_540 = 1.36e-11
+ mcrdlm2d_ca_w_1_120_s_3_500 = 1.94e-05  mcrdlm2d_cc_w_1_120_s_3_500 = 1.42e-11  mcrdlm2d_cf_w_1_120_s_3_500 = 2.42e-11
+ mcrdlm2p1_ca_w_0_140_s_0_140 = 2.15e-05  mcrdlm2p1_cc_w_0_140_s_0_140 = 8.78e-11  mcrdlm2p1_cf_w_0_140_s_0_140 = 1.83e-12
+ mcrdlm2p1_ca_w_0_140_s_0_175 = 2.15e-05  mcrdlm2p1_cc_w_0_140_s_0_175 = 8.63e-11  mcrdlm2p1_cf_w_0_140_s_0_175 = 2.20e-12
+ mcrdlm2p1_ca_w_0_140_s_0_210 = 2.15e-05  mcrdlm2p1_cc_w_0_140_s_0_210 = 8.35e-11  mcrdlm2p1_cf_w_0_140_s_0_210 = 2.58e-12
+ mcrdlm2p1_ca_w_0_140_s_0_280 = 2.15e-05  mcrdlm2p1_cc_w_0_140_s_0_280 = 7.60e-11  mcrdlm2p1_cf_w_0_140_s_0_280 = 3.31e-12
+ mcrdlm2p1_ca_w_0_140_s_0_350 = 2.15e-05  mcrdlm2p1_cc_w_0_140_s_0_350 = 6.71e-11  mcrdlm2p1_cf_w_0_140_s_0_350 = 4.04e-12
+ mcrdlm2p1_ca_w_0_140_s_0_420 = 2.15e-05  mcrdlm2p1_cc_w_0_140_s_0_420 = 5.99e-11  mcrdlm2p1_cf_w_0_140_s_0_420 = 4.79e-12
+ mcrdlm2p1_ca_w_0_140_s_0_560 = 2.15e-05  mcrdlm2p1_cc_w_0_140_s_0_560 = 4.97e-11  mcrdlm2p1_cf_w_0_140_s_0_560 = 6.18e-12
+ mcrdlm2p1_ca_w_0_140_s_0_840 = 2.15e-05  mcrdlm2p1_cc_w_0_140_s_0_840 = 3.78e-11  mcrdlm2p1_cf_w_0_140_s_0_840 = 8.81e-12
+ mcrdlm2p1_ca_w_0_140_s_1_540 = 2.15e-05  mcrdlm2p1_cc_w_0_140_s_1_540 = 2.35e-11  mcrdlm2p1_cf_w_0_140_s_1_540 = 1.45e-11
+ mcrdlm2p1_ca_w_0_140_s_3_500 = 2.15e-05  mcrdlm2p1_cc_w_0_140_s_3_500 = 9.33e-12  mcrdlm2p1_cf_w_0_140_s_3_500 = 2.41e-11
+ mcrdlm2p1_ca_w_1_120_s_0_140 = 2.15e-05  mcrdlm2p1_cc_w_1_120_s_0_140 = 1.14e-10  mcrdlm2p1_cf_w_1_120_s_0_140 = 1.87e-12
+ mcrdlm2p1_ca_w_1_120_s_0_175 = 2.15e-05  mcrdlm2p1_cc_w_1_120_s_0_175 = 1.12e-10  mcrdlm2p1_cf_w_1_120_s_0_175 = 2.25e-12
+ mcrdlm2p1_ca_w_1_120_s_0_210 = 2.15e-05  mcrdlm2p1_cc_w_1_120_s_0_210 = 1.07e-10  mcrdlm2p1_cf_w_1_120_s_0_210 = 2.62e-12
+ mcrdlm2p1_ca_w_1_120_s_0_280 = 2.15e-05  mcrdlm2p1_cc_w_1_120_s_0_280 = 9.58e-11  mcrdlm2p1_cf_w_1_120_s_0_280 = 3.36e-12
+ mcrdlm2p1_ca_w_1_120_s_0_350 = 2.15e-05  mcrdlm2p1_cc_w_1_120_s_0_350 = 8.58e-11  mcrdlm2p1_cf_w_1_120_s_0_350 = 4.10e-12
+ mcrdlm2p1_ca_w_1_120_s_0_420 = 2.15e-05  mcrdlm2p1_cc_w_1_120_s_0_420 = 7.69e-11  mcrdlm2p1_cf_w_1_120_s_0_420 = 4.82e-12
+ mcrdlm2p1_ca_w_1_120_s_0_560 = 2.15e-05  mcrdlm2p1_cc_w_1_120_s_0_560 = 6.43e-11  mcrdlm2p1_cf_w_1_120_s_0_560 = 6.23e-12
+ mcrdlm2p1_ca_w_1_120_s_0_840 = 2.15e-05  mcrdlm2p1_cc_w_1_120_s_0_840 = 4.91e-11  mcrdlm2p1_cf_w_1_120_s_0_840 = 8.92e-12
+ mcrdlm2p1_ca_w_1_120_s_1_540 = 2.15e-05  mcrdlm2p1_cc_w_1_120_s_1_540 = 3.13e-11  mcrdlm2p1_cf_w_1_120_s_1_540 = 1.49e-11
+ mcrdlm2p1_ca_w_1_120_s_3_500 = 2.15e-05  mcrdlm2p1_cc_w_1_120_s_3_500 = 1.32e-11  mcrdlm2p1_cf_w_1_120_s_3_500 = 2.59e-11
+ mcrdlm2l1_ca_w_0_140_s_0_140 = 3.12e-05  mcrdlm2l1_cc_w_0_140_s_0_140 = 8.67e-11  mcrdlm2l1_cf_w_0_140_s_0_140 = 2.62e-12
+ mcrdlm2l1_ca_w_0_140_s_0_175 = 3.12e-05  mcrdlm2l1_cc_w_0_140_s_0_175 = 8.52e-11  mcrdlm2l1_cf_w_0_140_s_0_175 = 3.16e-12
+ mcrdlm2l1_ca_w_0_140_s_0_210 = 3.12e-05  mcrdlm2l1_cc_w_0_140_s_0_210 = 8.21e-11  mcrdlm2l1_cf_w_0_140_s_0_210 = 3.71e-12
+ mcrdlm2l1_ca_w_0_140_s_0_280 = 3.12e-05  mcrdlm2l1_cc_w_0_140_s_0_280 = 7.43e-11  mcrdlm2l1_cf_w_0_140_s_0_280 = 4.76e-12
+ mcrdlm2l1_ca_w_0_140_s_0_350 = 3.12e-05  mcrdlm2l1_cc_w_0_140_s_0_350 = 6.54e-11  mcrdlm2l1_cf_w_0_140_s_0_350 = 5.79e-12
+ mcrdlm2l1_ca_w_0_140_s_0_420 = 3.12e-05  mcrdlm2l1_cc_w_0_140_s_0_420 = 5.79e-11  mcrdlm2l1_cf_w_0_140_s_0_420 = 6.84e-12
+ mcrdlm2l1_ca_w_0_140_s_0_560 = 3.12e-05  mcrdlm2l1_cc_w_0_140_s_0_560 = 4.73e-11  mcrdlm2l1_cf_w_0_140_s_0_560 = 8.78e-12
+ mcrdlm2l1_ca_w_0_140_s_0_840 = 3.12e-05  mcrdlm2l1_cc_w_0_140_s_0_840 = 3.50e-11  mcrdlm2l1_cf_w_0_140_s_0_840 = 1.24e-11
+ mcrdlm2l1_ca_w_0_140_s_1_540 = 3.12e-05  mcrdlm2l1_cc_w_0_140_s_1_540 = 2.03e-11  mcrdlm2l1_cf_w_0_140_s_1_540 = 1.97e-11
+ mcrdlm2l1_ca_w_0_140_s_3_500 = 3.12e-05  mcrdlm2l1_cc_w_0_140_s_3_500 = 6.85e-12  mcrdlm2l1_cf_w_0_140_s_3_500 = 3.00e-11
+ mcrdlm2l1_ca_w_1_120_s_0_140 = 3.12e-05  mcrdlm2l1_cc_w_1_120_s_0_140 = 1.11e-10  mcrdlm2l1_cf_w_1_120_s_0_140 = 2.65e-12
+ mcrdlm2l1_ca_w_1_120_s_0_175 = 3.12e-05  mcrdlm2l1_cc_w_1_120_s_0_175 = 1.08e-10  mcrdlm2l1_cf_w_1_120_s_0_175 = 3.20e-12
+ mcrdlm2l1_ca_w_1_120_s_0_210 = 3.12e-05  mcrdlm2l1_cc_w_1_120_s_0_210 = 1.04e-10  mcrdlm2l1_cf_w_1_120_s_0_210 = 3.73e-12
+ mcrdlm2l1_ca_w_1_120_s_0_280 = 3.12e-05  mcrdlm2l1_cc_w_1_120_s_0_280 = 9.20e-11  mcrdlm2l1_cf_w_1_120_s_0_280 = 4.79e-12
+ mcrdlm2l1_ca_w_1_120_s_0_350 = 3.12e-05  mcrdlm2l1_cc_w_1_120_s_0_350 = 8.21e-11  mcrdlm2l1_cf_w_1_120_s_0_350 = 5.84e-12
+ mcrdlm2l1_ca_w_1_120_s_0_420 = 3.12e-05  mcrdlm2l1_cc_w_1_120_s_0_420 = 7.31e-11  mcrdlm2l1_cf_w_1_120_s_0_420 = 6.85e-12
+ mcrdlm2l1_ca_w_1_120_s_0_560 = 3.12e-05  mcrdlm2l1_cc_w_1_120_s_0_560 = 6.02e-11  mcrdlm2l1_cf_w_1_120_s_0_560 = 8.83e-12
+ mcrdlm2l1_ca_w_1_120_s_0_840 = 3.12e-05  mcrdlm2l1_cc_w_1_120_s_0_840 = 4.51e-11  mcrdlm2l1_cf_w_1_120_s_0_840 = 1.25e-11
+ mcrdlm2l1_ca_w_1_120_s_1_540 = 3.12e-05  mcrdlm2l1_cc_w_1_120_s_1_540 = 2.72e-11  mcrdlm2l1_cf_w_1_120_s_1_540 = 2.02e-11
+ mcrdlm2l1_ca_w_1_120_s_3_500 = 3.12e-05  mcrdlm2l1_cc_w_1_120_s_3_500 = 1.02e-11  mcrdlm2l1_cf_w_1_120_s_3_500 = 3.23e-11
+ mcrdlm2m1_ca_w_0_140_s_0_140 = 8.30e-05  mcrdlm2m1_cc_w_0_140_s_0_140 = 8.16e-11  mcrdlm2m1_cf_w_0_140_s_0_140 = 6.66e-12
+ mcrdlm2m1_ca_w_0_140_s_0_175 = 8.30e-05  mcrdlm2m1_cc_w_0_140_s_0_175 = 7.98e-11  mcrdlm2m1_cf_w_0_140_s_0_175 = 8.12e-12
+ mcrdlm2m1_ca_w_0_140_s_0_210 = 8.30e-05  mcrdlm2m1_cc_w_0_140_s_0_210 = 7.63e-11  mcrdlm2m1_cf_w_0_140_s_0_210 = 9.50e-12
+ mcrdlm2m1_ca_w_0_140_s_0_280 = 8.30e-05  mcrdlm2m1_cc_w_0_140_s_0_280 = 6.75e-11  mcrdlm2m1_cf_w_0_140_s_0_280 = 1.21e-11
+ mcrdlm2m1_ca_w_0_140_s_0_350 = 8.30e-05  mcrdlm2m1_cc_w_0_140_s_0_350 = 5.78e-11  mcrdlm2m1_cf_w_0_140_s_0_350 = 1.46e-11
+ mcrdlm2m1_ca_w_0_140_s_0_420 = 8.30e-05  mcrdlm2m1_cc_w_0_140_s_0_420 = 4.96e-11  mcrdlm2m1_cf_w_0_140_s_0_420 = 1.70e-11
+ mcrdlm2m1_ca_w_0_140_s_0_560 = 8.30e-05  mcrdlm2m1_cc_w_0_140_s_0_560 = 3.88e-11  mcrdlm2m1_cf_w_0_140_s_0_560 = 2.12e-11
+ mcrdlm2m1_ca_w_0_140_s_0_840 = 8.30e-05  mcrdlm2m1_cc_w_0_140_s_0_840 = 2.60e-11  mcrdlm2m1_cf_w_0_140_s_0_840 = 2.82e-11
+ mcrdlm2m1_ca_w_0_140_s_1_540 = 8.30e-05  mcrdlm2m1_cc_w_0_140_s_1_540 = 1.22e-11  mcrdlm2m1_cf_w_0_140_s_1_540 = 3.87e-11
+ mcrdlm2m1_ca_w_0_140_s_3_500 = 8.30e-05  mcrdlm2m1_cc_w_0_140_s_3_500 = 3.10e-12  mcrdlm2m1_cf_w_0_140_s_3_500 = 4.74e-11
+ mcrdlm2m1_ca_w_1_120_s_0_140 = 8.30e-05  mcrdlm2m1_cc_w_1_120_s_0_140 = 1.00e-10  mcrdlm2m1_cf_w_1_120_s_0_140 = 6.69e-12
+ mcrdlm2m1_ca_w_1_120_s_0_175 = 8.30e-05  mcrdlm2m1_cc_w_1_120_s_0_175 = 9.73e-11  mcrdlm2m1_cf_w_1_120_s_0_175 = 8.12e-12
+ mcrdlm2m1_ca_w_1_120_s_0_210 = 8.30e-05  mcrdlm2m1_cc_w_1_120_s_0_210 = 9.22e-11  mcrdlm2m1_cf_w_1_120_s_0_210 = 9.50e-12
+ mcrdlm2m1_ca_w_1_120_s_0_280 = 8.30e-05  mcrdlm2m1_cc_w_1_120_s_0_280 = 8.13e-11  mcrdlm2m1_cf_w_1_120_s_0_280 = 1.21e-11
+ mcrdlm2m1_ca_w_1_120_s_0_350 = 8.30e-05  mcrdlm2m1_cc_w_1_120_s_0_350 = 7.10e-11  mcrdlm2m1_cf_w_1_120_s_0_350 = 1.46e-11
+ mcrdlm2m1_ca_w_1_120_s_0_420 = 8.30e-05  mcrdlm2m1_cc_w_1_120_s_0_420 = 6.23e-11  mcrdlm2m1_cf_w_1_120_s_0_420 = 1.70e-11
+ mcrdlm2m1_ca_w_1_120_s_0_560 = 8.30e-05  mcrdlm2m1_cc_w_1_120_s_0_560 = 4.94e-11  mcrdlm2m1_cf_w_1_120_s_0_560 = 2.13e-11
+ mcrdlm2m1_ca_w_1_120_s_0_840 = 8.30e-05  mcrdlm2m1_cc_w_1_120_s_0_840 = 3.47e-11  mcrdlm2m1_cf_w_1_120_s_0_840 = 2.84e-11
+ mcrdlm2m1_ca_w_1_120_s_1_540 = 8.30e-05  mcrdlm2m1_cc_w_1_120_s_1_540 = 1.84e-11  mcrdlm2m1_cf_w_1_120_s_1_540 = 3.98e-11
+ mcrdlm2m1_ca_w_1_120_s_3_500 = 8.30e-05  mcrdlm2m1_cc_w_1_120_s_3_500 = 5.68e-12  mcrdlm2m1_cf_w_1_120_s_3_500 = 5.13e-11
+ mcm4m3f_ca_w_0_300_s_0_300 = 6.78e-05  mcm4m3f_cc_w_0_300_s_0_300 = 8.04e-11  mcm4m3f_cf_w_0_300_s_0_300 = 1.03e-11
+ mcm4m3f_ca_w_0_300_s_0_360 = 6.78e-05  mcm4m3f_cc_w_0_300_s_0_360 = 7.39e-11  mcm4m3f_cf_w_0_300_s_0_360 = 1.20e-11
+ mcm4m3f_ca_w_0_300_s_0_450 = 6.78e-05  mcm4m3f_cc_w_0_300_s_0_450 = 6.56e-11  mcm4m3f_cf_w_0_300_s_0_450 = 1.45e-11
+ mcm4m3f_ca_w_0_300_s_0_600 = 6.78e-05  mcm4m3f_cc_w_0_300_s_0_600 = 5.43e-11  mcm4m3f_cf_w_0_300_s_0_600 = 1.83e-11
+ mcm4m3f_ca_w_0_300_s_0_800 = 6.78e-05  mcm4m3f_cc_w_0_300_s_0_800 = 4.29e-11  mcm4m3f_cf_w_0_300_s_0_800 = 2.28e-11
+ mcm4m3f_ca_w_0_300_s_1_000 = 6.78e-05  mcm4m3f_cc_w_0_300_s_1_000 = 3.41e-11  mcm4m3f_cf_w_0_300_s_1_000 = 2.68e-11
+ mcm4m3f_ca_w_0_300_s_1_200 = 6.78e-05  mcm4m3f_cc_w_0_300_s_1_200 = 2.77e-11  mcm4m3f_cf_w_0_300_s_1_200 = 3.02e-11
+ mcm4m3f_ca_w_0_300_s_2_100 = 6.78e-05  mcm4m3f_cc_w_0_300_s_2_100 = 1.21e-11  mcm4m3f_cf_w_0_300_s_2_100 = 4.09e-11
+ mcm4m3f_ca_w_0_300_s_3_300 = 6.78e-05  mcm4m3f_cc_w_0_300_s_3_300 = 4.75e-12  mcm4m3f_cf_w_0_300_s_3_300 = 4.72e-11
+ mcm4m3f_ca_w_0_300_s_9_000 = 6.78e-05  mcm4m3f_cc_w_0_300_s_9_000 = 1.50e-13  mcm4m3f_cf_w_0_300_s_9_000 = 5.17e-11
+ mcm4m3f_ca_w_2_400_s_0_300 = 6.78e-05  mcm4m3f_cc_w_2_400_s_0_300 = 9.00e-11  mcm4m3f_cf_w_2_400_s_0_300 = 1.04e-11
+ mcm4m3f_ca_w_2_400_s_0_360 = 6.78e-05  mcm4m3f_cc_w_2_400_s_0_360 = 8.32e-11  mcm4m3f_cf_w_2_400_s_0_360 = 1.21e-11
+ mcm4m3f_ca_w_2_400_s_0_450 = 6.78e-05  mcm4m3f_cc_w_2_400_s_0_450 = 7.40e-11  mcm4m3f_cf_w_2_400_s_0_450 = 1.46e-11
+ mcm4m3f_ca_w_2_400_s_0_600 = 6.78e-05  mcm4m3f_cc_w_2_400_s_0_600 = 6.16e-11  mcm4m3f_cf_w_2_400_s_0_600 = 1.84e-11
+ mcm4m3f_ca_w_2_400_s_0_800 = 6.78e-05  mcm4m3f_cc_w_2_400_s_0_800 = 4.87e-11  mcm4m3f_cf_w_2_400_s_0_800 = 2.30e-11
+ mcm4m3f_ca_w_2_400_s_1_000 = 6.78e-05  mcm4m3f_cc_w_2_400_s_1_000 = 3.92e-11  mcm4m3f_cf_w_2_400_s_1_000 = 2.70e-11
+ mcm4m3f_ca_w_2_400_s_1_200 = 6.78e-05  mcm4m3f_cc_w_2_400_s_1_200 = 3.20e-11  mcm4m3f_cf_w_2_400_s_1_200 = 3.06e-11
+ mcm4m3f_ca_w_2_400_s_2_100 = 6.78e-05  mcm4m3f_cc_w_2_400_s_2_100 = 1.48e-11  mcm4m3f_cf_w_2_400_s_2_100 = 4.18e-11
+ mcm4m3f_ca_w_2_400_s_3_300 = 6.78e-05  mcm4m3f_cc_w_2_400_s_3_300 = 6.14e-12  mcm4m3f_cf_w_2_400_s_3_300 = 4.91e-11
+ mcm4m3f_ca_w_2_400_s_9_000 = 6.78e-05  mcm4m3f_cc_w_2_400_s_9_000 = 1.40e-13  mcm4m3f_cf_w_2_400_s_9_000 = 5.48e-11
+ mcm4m3d_ca_w_0_300_s_0_300 = 6.92e-05  mcm4m3d_cc_w_0_300_s_0_300 = 8.01e-11  mcm4m3d_cf_w_0_300_s_0_300 = 1.06e-11
+ mcm4m3d_ca_w_0_300_s_0_360 = 6.92e-05  mcm4m3d_cc_w_0_300_s_0_360 = 7.35e-11  mcm4m3d_cf_w_0_300_s_0_360 = 1.23e-11
+ mcm4m3d_ca_w_0_300_s_0_450 = 6.92e-05  mcm4m3d_cc_w_0_300_s_0_450 = 6.53e-11  mcm4m3d_cf_w_0_300_s_0_450 = 1.48e-11
+ mcm4m3d_ca_w_0_300_s_0_600 = 6.92e-05  mcm4m3d_cc_w_0_300_s_0_600 = 5.39e-11  mcm4m3d_cf_w_0_300_s_0_600 = 1.87e-11
+ mcm4m3d_ca_w_0_300_s_0_800 = 6.92e-05  mcm4m3d_cc_w_0_300_s_0_800 = 4.23e-11  mcm4m3d_cf_w_0_300_s_0_800 = 2.33e-11
+ mcm4m3d_ca_w_0_300_s_1_000 = 6.92e-05  mcm4m3d_cc_w_0_300_s_1_000 = 3.34e-11  mcm4m3d_cf_w_0_300_s_1_000 = 2.74e-11
+ mcm4m3d_ca_w_0_300_s_1_200 = 6.92e-05  mcm4m3d_cc_w_0_300_s_1_200 = 2.70e-11  mcm4m3d_cf_w_0_300_s_1_200 = 3.09e-11
+ mcm4m3d_ca_w_0_300_s_2_100 = 6.92e-05  mcm4m3d_cc_w_0_300_s_2_100 = 1.15e-11  mcm4m3d_cf_w_0_300_s_2_100 = 4.17e-11
+ mcm4m3d_ca_w_0_300_s_3_300 = 6.92e-05  mcm4m3d_cc_w_0_300_s_3_300 = 4.28e-12  mcm4m3d_cf_w_0_300_s_3_300 = 4.79e-11
+ mcm4m3d_ca_w_0_300_s_9_000 = 6.92e-05  mcm4m3d_cc_w_0_300_s_9_000 = 1.15e-13  mcm4m3d_cf_w_0_300_s_9_000 = 5.20e-11
+ mcm4m3d_ca_w_2_400_s_0_300 = 6.92e-05  mcm4m3d_cc_w_2_400_s_0_300 = 8.89e-11  mcm4m3d_cf_w_2_400_s_0_300 = 1.07e-11
+ mcm4m3d_ca_w_2_400_s_0_360 = 6.92e-05  mcm4m3d_cc_w_2_400_s_0_360 = 8.20e-11  mcm4m3d_cf_w_2_400_s_0_360 = 1.24e-11
+ mcm4m3d_ca_w_2_400_s_0_450 = 6.92e-05  mcm4m3d_cc_w_2_400_s_0_450 = 7.29e-11  mcm4m3d_cf_w_2_400_s_0_450 = 1.49e-11
+ mcm4m3d_ca_w_2_400_s_0_600 = 6.92e-05  mcm4m3d_cc_w_2_400_s_0_600 = 6.04e-11  mcm4m3d_cf_w_2_400_s_0_600 = 1.88e-11
+ mcm4m3d_ca_w_2_400_s_0_800 = 6.92e-05  mcm4m3d_cc_w_2_400_s_0_800 = 4.75e-11  mcm4m3d_cf_w_2_400_s_0_800 = 2.35e-11
+ mcm4m3d_ca_w_2_400_s_1_000 = 6.92e-05  mcm4m3d_cc_w_2_400_s_1_000 = 3.80e-11  mcm4m3d_cf_w_2_400_s_1_000 = 2.77e-11
+ mcm4m3d_ca_w_2_400_s_1_200 = 6.92e-05  mcm4m3d_cc_w_2_400_s_1_200 = 3.08e-11  mcm4m3d_cf_w_2_400_s_1_200 = 3.13e-11
+ mcm4m3d_ca_w_2_400_s_2_100 = 6.92e-05  mcm4m3d_cc_w_2_400_s_2_100 = 1.38e-11  mcm4m3d_cf_w_2_400_s_2_100 = 4.26e-11
+ mcm4m3d_ca_w_2_400_s_3_300 = 6.92e-05  mcm4m3d_cc_w_2_400_s_3_300 = 5.31e-12  mcm4m3d_cf_w_2_400_s_3_300 = 4.98e-11
+ mcm4m3d_ca_w_2_400_s_9_000 = 6.92e-05  mcm4m3d_cc_w_2_400_s_9_000 = 1.25e-13  mcm4m3d_cf_w_2_400_s_9_000 = 5.48e-11
+ mcm4m3p1_ca_w_0_300_s_0_300 = 7.02e-05  mcm4m3p1_cc_w_0_300_s_0_300 = 7.96e-11  mcm4m3p1_cf_w_0_300_s_0_300 = 1.07e-11
+ mcm4m3p1_ca_w_0_300_s_0_360 = 7.02e-05  mcm4m3p1_cc_w_0_300_s_0_360 = 7.33e-11  mcm4m3p1_cf_w_0_300_s_0_360 = 1.25e-11
+ mcm4m3p1_ca_w_0_300_s_0_450 = 7.02e-05  mcm4m3p1_cc_w_0_300_s_0_450 = 6.49e-11  mcm4m3p1_cf_w_0_300_s_0_450 = 1.51e-11
+ mcm4m3p1_ca_w_0_300_s_0_600 = 7.02e-05  mcm4m3p1_cc_w_0_300_s_0_600 = 5.35e-11  mcm4m3p1_cf_w_0_300_s_0_600 = 1.90e-11
+ mcm4m3p1_ca_w_0_300_s_0_800 = 7.02e-05  mcm4m3p1_cc_w_0_300_s_0_800 = 4.19e-11  mcm4m3p1_cf_w_0_300_s_0_800 = 2.37e-11
+ mcm4m3p1_ca_w_0_300_s_1_000 = 7.02e-05  mcm4m3p1_cc_w_0_300_s_1_000 = 3.32e-11  mcm4m3p1_cf_w_0_300_s_1_000 = 2.78e-11
+ mcm4m3p1_ca_w_0_300_s_1_200 = 7.02e-05  mcm4m3p1_cc_w_0_300_s_1_200 = 2.65e-11  mcm4m3p1_cf_w_0_300_s_1_200 = 3.14e-11
+ mcm4m3p1_ca_w_0_300_s_2_100 = 7.02e-05  mcm4m3p1_cc_w_0_300_s_2_100 = 1.11e-11  mcm4m3p1_cf_w_0_300_s_2_100 = 4.21e-11
+ mcm4m3p1_ca_w_0_300_s_3_300 = 7.02e-05  mcm4m3p1_cc_w_0_300_s_3_300 = 4.00e-12  mcm4m3p1_cf_w_0_300_s_3_300 = 4.84e-11
+ mcm4m3p1_ca_w_0_300_s_9_000 = 7.02e-05  mcm4m3p1_cc_w_0_300_s_9_000 = 1.10e-13  mcm4m3p1_cf_w_0_300_s_9_000 = 5.21e-11
+ mcm4m3p1_ca_w_2_400_s_0_300 = 7.02e-05  mcm4m3p1_cc_w_2_400_s_0_300 = 8.81e-11  mcm4m3p1_cf_w_2_400_s_0_300 = 1.09e-11
+ mcm4m3p1_ca_w_2_400_s_0_360 = 7.02e-05  mcm4m3p1_cc_w_2_400_s_0_360 = 8.13e-11  mcm4m3p1_cf_w_2_400_s_0_360 = 1.26e-11
+ mcm4m3p1_ca_w_2_400_s_0_450 = 7.02e-05  mcm4m3p1_cc_w_2_400_s_0_450 = 7.21e-11  mcm4m3p1_cf_w_2_400_s_0_450 = 1.51e-11
+ mcm4m3p1_ca_w_2_400_s_0_600 = 7.02e-05  mcm4m3p1_cc_w_2_400_s_0_600 = 5.96e-11  mcm4m3p1_cf_w_2_400_s_0_600 = 1.91e-11
+ mcm4m3p1_ca_w_2_400_s_0_800 = 7.02e-05  mcm4m3p1_cc_w_2_400_s_0_800 = 4.67e-11  mcm4m3p1_cf_w_2_400_s_0_800 = 2.39e-11
+ mcm4m3p1_ca_w_2_400_s_1_000 = 7.02e-05  mcm4m3p1_cc_w_2_400_s_1_000 = 3.72e-11  mcm4m3p1_cf_w_2_400_s_1_000 = 2.82e-11
+ mcm4m3p1_ca_w_2_400_s_1_200 = 7.02e-05  mcm4m3p1_cc_w_2_400_s_1_200 = 3.01e-11  mcm4m3p1_cf_w_2_400_s_1_200 = 3.18e-11
+ mcm4m3p1_ca_w_2_400_s_2_100 = 7.02e-05  mcm4m3p1_cc_w_2_400_s_2_100 = 1.31e-11  mcm4m3p1_cf_w_2_400_s_2_100 = 4.32e-11
+ mcm4m3p1_ca_w_2_400_s_3_300 = 7.02e-05  mcm4m3p1_cc_w_2_400_s_3_300 = 4.92e-12  mcm4m3p1_cf_w_2_400_s_3_300 = 5.02e-11
+ mcm4m3p1_ca_w_2_400_s_9_000 = 7.02e-05  mcm4m3p1_cc_w_2_400_s_9_000 = 1.05e-13  mcm4m3p1_cf_w_2_400_s_9_000 = 5.49e-11
+ mcm4m3l1_ca_w_0_300_s_0_300 = 7.39e-05  mcm4m3l1_cc_w_0_300_s_0_300 = 7.89e-11  mcm4m3l1_cf_w_0_300_s_0_300 = 1.13e-11
+ mcm4m3l1_ca_w_0_300_s_0_360 = 7.39e-05  mcm4m3l1_cc_w_0_300_s_0_360 = 7.23e-11  mcm4m3l1_cf_w_0_300_s_0_360 = 1.32e-11
+ mcm4m3l1_ca_w_0_300_s_0_450 = 7.39e-05  mcm4m3l1_cc_w_0_300_s_0_450 = 6.40e-11  mcm4m3l1_cf_w_0_300_s_0_450 = 1.59e-11
+ mcm4m3l1_ca_w_0_300_s_0_600 = 7.39e-05  mcm4m3l1_cc_w_0_300_s_0_600 = 5.24e-11  mcm4m3l1_cf_w_0_300_s_0_600 = 2.01e-11
+ mcm4m3l1_ca_w_0_300_s_0_800 = 7.39e-05  mcm4m3l1_cc_w_0_300_s_0_800 = 4.05e-11  mcm4m3l1_cf_w_0_300_s_0_800 = 2.50e-11
+ mcm4m3l1_ca_w_0_300_s_1_000 = 7.39e-05  mcm4m3l1_cc_w_0_300_s_1_000 = 3.16e-11  mcm4m3l1_cf_w_0_300_s_1_000 = 2.94e-11
+ mcm4m3l1_ca_w_0_300_s_1_200 = 7.39e-05  mcm4m3l1_cc_w_0_300_s_1_200 = 2.51e-11  mcm4m3l1_cf_w_0_300_s_1_200 = 3.31e-11
+ mcm4m3l1_ca_w_0_300_s_2_100 = 7.39e-05  mcm4m3l1_cc_w_0_300_s_2_100 = 9.72e-12  mcm4m3l1_cf_w_0_300_s_2_100 = 4.40e-11
+ mcm4m3l1_ca_w_0_300_s_3_300 = 7.39e-05  mcm4m3l1_cc_w_0_300_s_3_300 = 3.13e-12  mcm4m3l1_cf_w_0_300_s_3_300 = 5.00e-11
+ mcm4m3l1_ca_w_0_300_s_9_000 = 7.39e-05  mcm4m3l1_cc_w_0_300_s_9_000 = 4.50e-14  mcm4m3l1_cf_w_0_300_s_9_000 = 5.30e-11
+ mcm4m3l1_ca_w_2_400_s_0_300 = 7.39e-05  mcm4m3l1_cc_w_2_400_s_0_300 = 8.56e-11  mcm4m3l1_cf_w_2_400_s_0_300 = 1.15e-11
+ mcm4m3l1_ca_w_2_400_s_0_360 = 7.39e-05  mcm4m3l1_cc_w_2_400_s_0_360 = 7.88e-11  mcm4m3l1_cf_w_2_400_s_0_360 = 1.33e-11
+ mcm4m3l1_ca_w_2_400_s_0_450 = 7.39e-05  mcm4m3l1_cc_w_2_400_s_0_450 = 6.96e-11  mcm4m3l1_cf_w_2_400_s_0_450 = 1.60e-11
+ mcm4m3l1_ca_w_2_400_s_0_600 = 7.39e-05  mcm4m3l1_cc_w_2_400_s_0_600 = 5.70e-11  mcm4m3l1_cf_w_2_400_s_0_600 = 2.02e-11
+ mcm4m3l1_ca_w_2_400_s_0_800 = 7.39e-05  mcm4m3l1_cc_w_2_400_s_0_800 = 4.41e-11  mcm4m3l1_cf_w_2_400_s_0_800 = 2.52e-11
+ mcm4m3l1_ca_w_2_400_s_1_000 = 7.39e-05  mcm4m3l1_cc_w_2_400_s_1_000 = 3.46e-11  mcm4m3l1_cf_w_2_400_s_1_000 = 2.97e-11
+ mcm4m3l1_ca_w_2_400_s_1_200 = 7.39e-05  mcm4m3l1_cc_w_2_400_s_1_200 = 2.75e-11  mcm4m3l1_cf_w_2_400_s_1_200 = 3.35e-11
+ mcm4m3l1_ca_w_2_400_s_2_100 = 7.39e-05  mcm4m3l1_cc_w_2_400_s_2_100 = 1.10e-11  mcm4m3l1_cf_w_2_400_s_2_100 = 4.50e-11
+ mcm4m3l1_ca_w_2_400_s_3_300 = 7.39e-05  mcm4m3l1_cc_w_2_400_s_3_300 = 3.59e-12  mcm4m3l1_cf_w_2_400_s_3_300 = 5.16e-11
+ mcm4m3l1_ca_w_2_400_s_9_000 = 7.39e-05  mcm4m3l1_cc_w_2_400_s_9_000 = 7.00e-14  mcm4m3l1_cf_w_2_400_s_9_000 = 5.51e-11
+ mcm4m3m1_ca_w_0_300_s_0_300 = 8.33e-05  mcm4m3m1_cc_w_0_300_s_0_300 = 7.67e-11  mcm4m3m1_cf_w_0_300_s_0_300 = 1.29e-11
+ mcm4m3m1_ca_w_0_300_s_0_360 = 8.33e-05  mcm4m3m1_cc_w_0_300_s_0_360 = 6.99e-11  mcm4m3m1_cf_w_0_300_s_0_360 = 1.50e-11
+ mcm4m3m1_ca_w_0_300_s_0_450 = 8.33e-05  mcm4m3m1_cc_w_0_300_s_0_450 = 6.15e-11  mcm4m3m1_cf_w_0_300_s_0_450 = 1.80e-11
+ mcm4m3m1_ca_w_0_300_s_0_600 = 8.33e-05  mcm4m3m1_cc_w_0_300_s_0_600 = 4.94e-11  mcm4m3m1_cf_w_0_300_s_0_600 = 2.27e-11
+ mcm4m3m1_ca_w_0_300_s_0_800 = 8.33e-05  mcm4m3m1_cc_w_0_300_s_0_800 = 3.73e-11  mcm4m3m1_cf_w_0_300_s_0_800 = 2.82e-11
+ mcm4m3m1_ca_w_0_300_s_1_000 = 8.33e-05  mcm4m3m1_cc_w_0_300_s_1_000 = 2.84e-11  mcm4m3m1_cf_w_0_300_s_1_000 = 3.31e-11
+ mcm4m3m1_ca_w_0_300_s_1_200 = 8.33e-05  mcm4m3m1_cc_w_0_300_s_1_200 = 2.19e-11  mcm4m3m1_cf_w_0_300_s_1_200 = 3.72e-11
+ mcm4m3m1_ca_w_0_300_s_2_100 = 8.33e-05  mcm4m3m1_cc_w_0_300_s_2_100 = 7.24e-12  mcm4m3m1_cf_w_0_300_s_2_100 = 4.83e-11
+ mcm4m3m1_ca_w_0_300_s_3_300 = 8.33e-05  mcm4m3m1_cc_w_0_300_s_3_300 = 1.77e-12  mcm4m3m1_cf_w_0_300_s_3_300 = 5.33e-11
+ mcm4m3m1_ca_w_0_300_s_9_000 = 8.33e-05  mcm4m3m1_cc_w_0_300_s_9_000 = 2.50e-14  mcm4m3m1_cf_w_0_300_s_9_000 = 5.52e-11
+ mcm4m3m1_ca_w_2_400_s_0_300 = 8.33e-05  mcm4m3m1_cc_w_2_400_s_0_300 = 8.08e-11  mcm4m3m1_cf_w_2_400_s_0_300 = 1.30e-11
+ mcm4m3m1_ca_w_2_400_s_0_360 = 8.33e-05  mcm4m3m1_cc_w_2_400_s_0_360 = 7.39e-11  mcm4m3m1_cf_w_2_400_s_0_360 = 1.51e-11
+ mcm4m3m1_ca_w_2_400_s_0_450 = 8.33e-05  mcm4m3m1_cc_w_2_400_s_0_450 = 6.47e-11  mcm4m3m1_cf_w_2_400_s_0_450 = 1.81e-11
+ mcm4m3m1_ca_w_2_400_s_0_600 = 8.33e-05  mcm4m3m1_cc_w_2_400_s_0_600 = 5.22e-11  mcm4m3m1_cf_w_2_400_s_0_600 = 2.29e-11
+ mcm4m3m1_ca_w_2_400_s_0_800 = 8.33e-05  mcm4m3m1_cc_w_2_400_s_0_800 = 3.94e-11  mcm4m3m1_cf_w_2_400_s_0_800 = 2.85e-11
+ mcm4m3m1_ca_w_2_400_s_1_000 = 8.33e-05  mcm4m3m1_cc_w_2_400_s_1_000 = 3.00e-11  mcm4m3m1_cf_w_2_400_s_1_000 = 3.34e-11
+ mcm4m3m1_ca_w_2_400_s_1_200 = 8.33e-05  mcm4m3m1_cc_w_2_400_s_1_200 = 2.31e-11  mcm4m3m1_cf_w_2_400_s_1_200 = 3.76e-11
+ mcm4m3m1_ca_w_2_400_s_2_100 = 8.33e-05  mcm4m3m1_cc_w_2_400_s_2_100 = 7.71e-12  mcm4m3m1_cf_w_2_400_s_2_100 = 4.91e-11
+ mcm4m3m1_ca_w_2_400_s_3_300 = 8.33e-05  mcm4m3m1_cc_w_2_400_s_3_300 = 1.90e-12  mcm4m3m1_cf_w_2_400_s_3_300 = 5.46e-11
+ mcm4m3m1_ca_w_2_400_s_9_000 = 8.33e-05  mcm4m3m1_cc_w_2_400_s_9_000 = 0.00e+00  mcm4m3m1_cf_w_2_400_s_9_000 = 5.65e-11
+ mcm4m3m2_ca_w_0_300_s_0_300 = 1.17e-04  mcm4m3m2_cc_w_0_300_s_0_300 = 7.03e-11  mcm4m3m2_cf_w_0_300_s_0_300 = 1.80e-11
+ mcm4m3m2_ca_w_0_300_s_0_360 = 1.17e-04  mcm4m3m2_cc_w_0_300_s_0_360 = 6.36e-11  mcm4m3m2_cf_w_0_300_s_0_360 = 2.09e-11
+ mcm4m3m2_ca_w_0_300_s_0_450 = 1.17e-04  mcm4m3m2_cc_w_0_300_s_0_450 = 5.47e-11  mcm4m3m2_cf_w_0_300_s_0_450 = 2.49e-11
+ mcm4m3m2_ca_w_0_300_s_0_600 = 1.17e-04  mcm4m3m2_cc_w_0_300_s_0_600 = 4.25e-11  mcm4m3m2_cf_w_0_300_s_0_600 = 3.11e-11
+ mcm4m3m2_ca_w_0_300_s_0_800 = 1.17e-04  mcm4m3m2_cc_w_0_300_s_0_800 = 3.04e-11  mcm4m3m2_cf_w_0_300_s_0_800 = 3.81e-11
+ mcm4m3m2_ca_w_0_300_s_1_000 = 1.17e-04  mcm4m3m2_cc_w_0_300_s_1_000 = 2.16e-11  mcm4m3m2_cf_w_0_300_s_1_000 = 4.40e-11
+ mcm4m3m2_ca_w_0_300_s_1_200 = 1.17e-04  mcm4m3m2_cc_w_0_300_s_1_200 = 1.55e-11  mcm4m3m2_cf_w_0_300_s_1_200 = 4.85e-11
+ mcm4m3m2_ca_w_0_300_s_2_100 = 1.17e-04  mcm4m3m2_cc_w_0_300_s_2_100 = 3.63e-12  mcm4m3m2_cf_w_0_300_s_2_100 = 5.87e-11
+ mcm4m3m2_ca_w_0_300_s_3_300 = 1.17e-04  mcm4m3m2_cc_w_0_300_s_3_300 = 6.05e-13  mcm4m3m2_cf_w_0_300_s_3_300 = 6.19e-11
+ mcm4m3m2_ca_w_0_300_s_9_000 = 1.17e-04  mcm4m3m2_cc_w_0_300_s_9_000 = 3.50e-14  mcm4m3m2_cf_w_0_300_s_9_000 = 6.23e-11
+ mcm4m3m2_ca_w_2_400_s_0_300 = 1.17e-04  mcm4m3m2_cc_w_2_400_s_0_300 = 7.16e-11  mcm4m3m2_cf_w_2_400_s_0_300 = 1.81e-11
+ mcm4m3m2_ca_w_2_400_s_0_360 = 1.17e-04  mcm4m3m2_cc_w_2_400_s_0_360 = 6.49e-11  mcm4m3m2_cf_w_2_400_s_0_360 = 2.10e-11
+ mcm4m3m2_ca_w_2_400_s_0_450 = 1.17e-04  mcm4m3m2_cc_w_2_400_s_0_450 = 5.58e-11  mcm4m3m2_cf_w_2_400_s_0_450 = 2.50e-11
+ mcm4m3m2_ca_w_2_400_s_0_600 = 1.17e-04  mcm4m3m2_cc_w_2_400_s_0_600 = 4.34e-11  mcm4m3m2_cf_w_2_400_s_0_600 = 3.12e-11
+ mcm4m3m2_ca_w_2_400_s_0_800 = 1.17e-04  mcm4m3m2_cc_w_2_400_s_0_800 = 3.10e-11  mcm4m3m2_cf_w_2_400_s_0_800 = 3.84e-11
+ mcm4m3m2_ca_w_2_400_s_1_000 = 1.17e-04  mcm4m3m2_cc_w_2_400_s_1_000 = 2.22e-11  mcm4m3m2_cf_w_2_400_s_1_000 = 4.44e-11
+ mcm4m3m2_ca_w_2_400_s_1_200 = 1.17e-04  mcm4m3m2_cc_w_2_400_s_1_200 = 1.59e-11  mcm4m3m2_cf_w_2_400_s_1_200 = 4.90e-11
+ mcm4m3m2_ca_w_2_400_s_2_100 = 1.17e-04  mcm4m3m2_cc_w_2_400_s_2_100 = 3.65e-12  mcm4m3m2_cf_w_2_400_s_2_100 = 5.95e-11
+ mcm4m3m2_ca_w_2_400_s_3_300 = 1.17e-04  mcm4m3m2_cc_w_2_400_s_3_300 = 6.00e-13  mcm4m3m2_cf_w_2_400_s_3_300 = 6.24e-11
+ mcm4m3m2_ca_w_2_400_s_9_000 = 1.17e-04  mcm4m3m2_cc_w_2_400_s_9_000 = 0.00e+00  mcm4m3m2_cf_w_2_400_s_9_000 = 6.29e-11
+ mcm5m3f_ca_w_0_300_s_0_300 = 2.69e-05  mcm5m3f_cc_w_0_300_s_0_300 = 8.78e-11  mcm5m3f_cf_w_0_300_s_0_300 = 4.51e-12
+ mcm5m3f_ca_w_0_300_s_0_360 = 2.69e-05  mcm5m3f_cc_w_0_300_s_0_360 = 8.19e-11  mcm5m3f_cf_w_0_300_s_0_360 = 5.28e-12
+ mcm5m3f_ca_w_0_300_s_0_450 = 2.69e-05  mcm5m3f_cc_w_0_300_s_0_450 = 7.41e-11  mcm5m3f_cf_w_0_300_s_0_450 = 6.47e-12
+ mcm5m3f_ca_w_0_300_s_0_600 = 2.69e-05  mcm5m3f_cc_w_0_300_s_0_600 = 6.34e-11  mcm5m3f_cf_w_0_300_s_0_600 = 8.36e-12
+ mcm5m3f_ca_w_0_300_s_0_800 = 2.69e-05  mcm5m3f_cc_w_0_300_s_0_800 = 5.26e-11  mcm5m3f_cf_w_0_300_s_0_800 = 1.06e-11
+ mcm5m3f_ca_w_0_300_s_1_000 = 2.69e-05  mcm5m3f_cc_w_0_300_s_1_000 = 4.40e-11  mcm5m3f_cf_w_0_300_s_1_000 = 1.29e-11
+ mcm5m3f_ca_w_0_300_s_1_200 = 2.69e-05  mcm5m3f_cc_w_0_300_s_1_200 = 3.75e-11  mcm5m3f_cf_w_0_300_s_1_200 = 1.50e-11
+ mcm5m3f_ca_w_0_300_s_2_100 = 2.69e-05  mcm5m3f_cc_w_0_300_s_2_100 = 2.06e-11  mcm5m3f_cf_w_0_300_s_2_100 = 2.31e-11
+ mcm5m3f_ca_w_0_300_s_3_300 = 2.69e-05  mcm5m3f_cc_w_0_300_s_3_300 = 1.04e-11  mcm5m3f_cf_w_0_300_s_3_300 = 3.00e-11
+ mcm5m3f_ca_w_0_300_s_9_000 = 2.69e-05  mcm5m3f_cc_w_0_300_s_9_000 = 5.80e-13  mcm5m3f_cf_w_0_300_s_9_000 = 3.87e-11
+ mcm5m3f_ca_w_2_400_s_0_300 = 2.69e-05  mcm5m3f_cc_w_2_400_s_0_300 = 1.03e-10  mcm5m3f_cf_w_2_400_s_0_300 = 4.55e-12
+ mcm5m3f_ca_w_2_400_s_0_360 = 2.69e-05  mcm5m3f_cc_w_2_400_s_0_360 = 9.63e-11  mcm5m3f_cf_w_2_400_s_0_360 = 5.33e-12
+ mcm5m3f_ca_w_2_400_s_0_450 = 2.69e-05  mcm5m3f_cc_w_2_400_s_0_450 = 8.71e-11  mcm5m3f_cf_w_2_400_s_0_450 = 6.47e-12
+ mcm5m3f_ca_w_2_400_s_0_600 = 2.69e-05  mcm5m3f_cc_w_2_400_s_0_600 = 7.44e-11  mcm5m3f_cf_w_2_400_s_0_600 = 8.32e-12
+ mcm5m3f_ca_w_2_400_s_0_800 = 2.69e-05  mcm5m3f_cc_w_2_400_s_0_800 = 6.16e-11  mcm5m3f_cf_w_2_400_s_0_800 = 1.07e-11
+ mcm5m3f_ca_w_2_400_s_1_000 = 2.69e-05  mcm5m3f_cc_w_2_400_s_1_000 = 5.16e-11  mcm5m3f_cf_w_2_400_s_1_000 = 1.30e-11
+ mcm5m3f_ca_w_2_400_s_1_200 = 2.69e-05  mcm5m3f_cc_w_2_400_s_1_200 = 4.40e-11  mcm5m3f_cf_w_2_400_s_1_200 = 1.52e-11
+ mcm5m3f_ca_w_2_400_s_2_100 = 2.69e-05  mcm5m3f_cc_w_2_400_s_2_100 = 2.45e-11  mcm5m3f_cf_w_2_400_s_2_100 = 2.36e-11
+ mcm5m3f_ca_w_2_400_s_3_300 = 2.69e-05  mcm5m3f_cc_w_2_400_s_3_300 = 1.26e-11  mcm5m3f_cf_w_2_400_s_3_300 = 3.15e-11
+ mcm5m3f_ca_w_2_400_s_9_000 = 2.69e-05  mcm5m3f_cc_w_2_400_s_9_000 = 7.30e-13  mcm5m3f_cf_w_2_400_s_9_000 = 4.19e-11
+ mcm5m3d_ca_w_0_300_s_0_300 = 2.83e-05  mcm5m3d_cc_w_0_300_s_0_300 = 8.74e-11  mcm5m3d_cf_w_0_300_s_0_300 = 4.75e-12
+ mcm5m3d_ca_w_0_300_s_0_360 = 2.83e-05  mcm5m3d_cc_w_0_300_s_0_360 = 8.16e-11  mcm5m3d_cf_w_0_300_s_0_360 = 5.57e-12
+ mcm5m3d_ca_w_0_300_s_0_450 = 2.83e-05  mcm5m3d_cc_w_0_300_s_0_450 = 7.37e-11  mcm5m3d_cf_w_0_300_s_0_450 = 6.81e-12
+ mcm5m3d_ca_w_0_300_s_0_600 = 2.83e-05  mcm5m3d_cc_w_0_300_s_0_600 = 6.29e-11  mcm5m3d_cf_w_0_300_s_0_600 = 8.79e-12
+ mcm5m3d_ca_w_0_300_s_0_800 = 2.83e-05  mcm5m3d_cc_w_0_300_s_0_800 = 5.20e-11  mcm5m3d_cf_w_0_300_s_0_800 = 1.12e-11
+ mcm5m3d_ca_w_0_300_s_1_000 = 2.83e-05  mcm5m3d_cc_w_0_300_s_1_000 = 4.33e-11  mcm5m3d_cf_w_0_300_s_1_000 = 1.35e-11
+ mcm5m3d_ca_w_0_300_s_1_200 = 2.83e-05  mcm5m3d_cc_w_0_300_s_1_200 = 3.68e-11  mcm5m3d_cf_w_0_300_s_1_200 = 1.58e-11
+ mcm5m3d_ca_w_0_300_s_2_100 = 2.83e-05  mcm5m3d_cc_w_0_300_s_2_100 = 1.98e-11  mcm5m3d_cf_w_0_300_s_2_100 = 2.41e-11
+ mcm5m3d_ca_w_0_300_s_3_300 = 2.83e-05  mcm5m3d_cc_w_0_300_s_3_300 = 9.70e-12  mcm5m3d_cf_w_0_300_s_3_300 = 3.11e-11
+ mcm5m3d_ca_w_0_300_s_9_000 = 2.83e-05  mcm5m3d_cc_w_0_300_s_9_000 = 4.55e-13  mcm5m3d_cf_w_0_300_s_9_000 = 3.93e-11
+ mcm5m3d_ca_w_2_400_s_0_300 = 2.83e-05  mcm5m3d_cc_w_2_400_s_0_300 = 1.02e-10  mcm5m3d_cf_w_2_400_s_0_300 = 4.80e-12
+ mcm5m3d_ca_w_2_400_s_0_360 = 2.83e-05  mcm5m3d_cc_w_2_400_s_0_360 = 9.51e-11  mcm5m3d_cf_w_2_400_s_0_360 = 5.62e-12
+ mcm5m3d_ca_w_2_400_s_0_450 = 2.83e-05  mcm5m3d_cc_w_2_400_s_0_450 = 8.59e-11  mcm5m3d_cf_w_2_400_s_0_450 = 6.81e-12
+ mcm5m3d_ca_w_2_400_s_0_600 = 2.83e-05  mcm5m3d_cc_w_2_400_s_0_600 = 7.32e-11  mcm5m3d_cf_w_2_400_s_0_600 = 8.76e-12
+ mcm5m3d_ca_w_2_400_s_0_800 = 2.83e-05  mcm5m3d_cc_w_2_400_s_0_800 = 6.03e-11  mcm5m3d_cf_w_2_400_s_0_800 = 1.13e-11
+ mcm5m3d_ca_w_2_400_s_1_000 = 2.83e-05  mcm5m3d_cc_w_2_400_s_1_000 = 5.04e-11  mcm5m3d_cf_w_2_400_s_1_000 = 1.37e-11
+ mcm5m3d_ca_w_2_400_s_1_200 = 2.83e-05  mcm5m3d_cc_w_2_400_s_1_200 = 4.28e-11  mcm5m3d_cf_w_2_400_s_1_200 = 1.60e-11
+ mcm5m3d_ca_w_2_400_s_2_100 = 2.83e-05  mcm5m3d_cc_w_2_400_s_2_100 = 2.33e-11  mcm5m3d_cf_w_2_400_s_2_100 = 2.47e-11
+ mcm5m3d_ca_w_2_400_s_3_300 = 2.83e-05  mcm5m3d_cc_w_2_400_s_3_300 = 1.16e-11  mcm5m3d_cf_w_2_400_s_3_300 = 3.26e-11
+ mcm5m3d_ca_w_2_400_s_9_000 = 2.83e-05  mcm5m3d_cc_w_2_400_s_9_000 = 5.60e-13  mcm5m3d_cf_w_2_400_s_9_000 = 4.24e-11
+ mcm5m3p1_ca_w_0_300_s_0_300 = 2.93e-05  mcm5m3p1_cc_w_0_300_s_0_300 = 8.71e-11  mcm5m3p1_cf_w_0_300_s_0_300 = 4.92e-12
+ mcm5m3p1_ca_w_0_300_s_0_360 = 2.93e-05  mcm5m3p1_cc_w_0_300_s_0_360 = 8.13e-11  mcm5m3p1_cf_w_0_300_s_0_360 = 5.76e-12
+ mcm5m3p1_ca_w_0_300_s_0_450 = 2.93e-05  mcm5m3p1_cc_w_0_300_s_0_450 = 7.34e-11  mcm5m3p1_cf_w_0_300_s_0_450 = 7.04e-12
+ mcm5m3p1_ca_w_0_300_s_0_600 = 2.93e-05  mcm5m3p1_cc_w_0_300_s_0_600 = 6.25e-11  mcm5m3p1_cf_w_0_300_s_0_600 = 9.09e-12
+ mcm5m3p1_ca_w_0_300_s_0_800 = 2.93e-05  mcm5m3p1_cc_w_0_300_s_0_800 = 5.16e-11  mcm5m3p1_cf_w_0_300_s_0_800 = 1.16e-11
+ mcm5m3p1_ca_w_0_300_s_1_000 = 2.93e-05  mcm5m3p1_cc_w_0_300_s_1_000 = 4.29e-11  mcm5m3p1_cf_w_0_300_s_1_000 = 1.40e-11
+ mcm5m3p1_ca_w_0_300_s_1_200 = 2.93e-05  mcm5m3p1_cc_w_0_300_s_1_200 = 3.63e-11  mcm5m3p1_cf_w_0_300_s_1_200 = 1.63e-11
+ mcm5m3p1_ca_w_0_300_s_2_100 = 2.93e-05  mcm5m3p1_cc_w_0_300_s_2_100 = 1.92e-11  mcm5m3p1_cf_w_0_300_s_2_100 = 2.47e-11
+ mcm5m3p1_ca_w_0_300_s_3_300 = 2.93e-05  mcm5m3p1_cc_w_0_300_s_3_300 = 9.24e-12  mcm5m3p1_cf_w_0_300_s_3_300 = 3.19e-11
+ mcm5m3p1_ca_w_0_300_s_9_000 = 2.93e-05  mcm5m3p1_cc_w_0_300_s_9_000 = 3.90e-13  mcm5m3p1_cf_w_0_300_s_9_000 = 3.97e-11
+ mcm5m3p1_ca_w_2_400_s_0_300 = 2.93e-05  mcm5m3p1_cc_w_2_400_s_0_300 = 1.02e-10  mcm5m3p1_cf_w_2_400_s_0_300 = 4.99e-12
+ mcm5m3p1_ca_w_2_400_s_0_360 = 2.93e-05  mcm5m3p1_cc_w_2_400_s_0_360 = 9.43e-11  mcm5m3p1_cf_w_2_400_s_0_360 = 5.84e-12
+ mcm5m3p1_ca_w_2_400_s_0_450 = 2.93e-05  mcm5m3p1_cc_w_2_400_s_0_450 = 8.52e-11  mcm5m3p1_cf_w_2_400_s_0_450 = 7.07e-12
+ mcm5m3p1_ca_w_2_400_s_0_600 = 2.93e-05  mcm5m3p1_cc_w_2_400_s_0_600 = 7.24e-11  mcm5m3p1_cf_w_2_400_s_0_600 = 9.08e-12
+ mcm5m3p1_ca_w_2_400_s_0_800 = 2.93e-05  mcm5m3p1_cc_w_2_400_s_0_800 = 5.95e-11  mcm5m3p1_cf_w_2_400_s_0_800 = 1.17e-11
+ mcm5m3p1_ca_w_2_400_s_1_000 = 2.93e-05  mcm5m3p1_cc_w_2_400_s_1_000 = 4.95e-11  mcm5m3p1_cf_w_2_400_s_1_000 = 1.42e-11
+ mcm5m3p1_ca_w_2_400_s_1_200 = 2.93e-05  mcm5m3p1_cc_w_2_400_s_1_200 = 4.20e-11  mcm5m3p1_cf_w_2_400_s_1_200 = 1.66e-11
+ mcm5m3p1_ca_w_2_400_s_2_100 = 2.93e-05  mcm5m3p1_cc_w_2_400_s_2_100 = 2.25e-11  mcm5m3p1_cf_w_2_400_s_2_100 = 2.55e-11
+ mcm5m3p1_ca_w_2_400_s_3_300 = 2.93e-05  mcm5m3p1_cc_w_2_400_s_3_300 = 1.09e-11  mcm5m3p1_cf_w_2_400_s_3_300 = 3.34e-11
+ mcm5m3p1_ca_w_2_400_s_9_000 = 2.93e-05  mcm5m3p1_cc_w_2_400_s_9_000 = 4.50e-13  mcm5m3p1_cf_w_2_400_s_9_000 = 4.28e-11
+ mcm5m3l1_ca_w_0_300_s_0_300 = 3.30e-05  mcm5m3l1_cc_w_0_300_s_0_300 = 8.62e-11  mcm5m3l1_cf_w_0_300_s_0_300 = 5.53e-12
+ mcm5m3l1_ca_w_0_300_s_0_360 = 3.30e-05  mcm5m3l1_cc_w_0_300_s_0_360 = 8.03e-11  mcm5m3l1_cf_w_0_300_s_0_360 = 6.47e-12
+ mcm5m3l1_ca_w_0_300_s_0_450 = 3.30e-05  mcm5m3l1_cc_w_0_300_s_0_450 = 7.23e-11  mcm5m3l1_cf_w_0_300_s_0_450 = 7.90e-12
+ mcm5m3l1_ca_w_0_300_s_0_600 = 3.30e-05  mcm5m3l1_cc_w_0_300_s_0_600 = 6.13e-11  mcm5m3l1_cf_w_0_300_s_0_600 = 1.02e-11
+ mcm5m3l1_ca_w_0_300_s_0_800 = 3.30e-05  mcm5m3l1_cc_w_0_300_s_0_800 = 5.02e-11  mcm5m3l1_cf_w_0_300_s_0_800 = 1.29e-11
+ mcm5m3l1_ca_w_0_300_s_1_000 = 3.30e-05  mcm5m3l1_cc_w_0_300_s_1_000 = 4.14e-11  mcm5m3l1_cf_w_0_300_s_1_000 = 1.56e-11
+ mcm5m3l1_ca_w_0_300_s_1_200 = 3.30e-05  mcm5m3l1_cc_w_0_300_s_1_200 = 3.47e-11  mcm5m3l1_cf_w_0_300_s_1_200 = 1.81e-11
+ mcm5m3l1_ca_w_0_300_s_2_100 = 3.30e-05  mcm5m3l1_cc_w_0_300_s_2_100 = 1.75e-11  mcm5m3l1_cf_w_0_300_s_2_100 = 2.72e-11
+ mcm5m3l1_ca_w_0_300_s_3_300 = 3.30e-05  mcm5m3l1_cc_w_0_300_s_3_300 = 7.85e-12  mcm5m3l1_cf_w_0_300_s_3_300 = 3.44e-11
+ mcm5m3l1_ca_w_0_300_s_9_000 = 3.30e-05  mcm5m3l1_cc_w_0_300_s_9_000 = 2.45e-13  mcm5m3l1_cf_w_0_300_s_9_000 = 4.14e-11
+ mcm5m3l1_ca_w_2_400_s_0_300 = 3.30e-05  mcm5m3l1_cc_w_2_400_s_0_300 = 9.89e-11  mcm5m3l1_cf_w_2_400_s_0_300 = 5.58e-12
+ mcm5m3l1_ca_w_2_400_s_0_360 = 3.30e-05  mcm5m3l1_cc_w_2_400_s_0_360 = 9.18e-11  mcm5m3l1_cf_w_2_400_s_0_360 = 6.53e-12
+ mcm5m3l1_ca_w_2_400_s_0_450 = 3.30e-05  mcm5m3l1_cc_w_2_400_s_0_450 = 8.26e-11  mcm5m3l1_cf_w_2_400_s_0_450 = 7.91e-12
+ mcm5m3l1_ca_w_2_400_s_0_600 = 3.30e-05  mcm5m3l1_cc_w_2_400_s_0_600 = 6.98e-11  mcm5m3l1_cf_w_2_400_s_0_600 = 1.02e-11
+ mcm5m3l1_ca_w_2_400_s_0_800 = 3.30e-05  mcm5m3l1_cc_w_2_400_s_0_800 = 5.69e-11  mcm5m3l1_cf_w_2_400_s_0_800 = 1.30e-11
+ mcm5m3l1_ca_w_2_400_s_1_000 = 3.30e-05  mcm5m3l1_cc_w_2_400_s_1_000 = 4.69e-11  mcm5m3l1_cf_w_2_400_s_1_000 = 1.58e-11
+ mcm5m3l1_ca_w_2_400_s_1_200 = 3.30e-05  mcm5m3l1_cc_w_2_400_s_1_200 = 3.94e-11  mcm5m3l1_cf_w_2_400_s_1_200 = 1.84e-11
+ mcm5m3l1_ca_w_2_400_s_2_100 = 3.30e-05  mcm5m3l1_cc_w_2_400_s_2_100 = 2.01e-11  mcm5m3l1_cf_w_2_400_s_2_100 = 2.79e-11
+ mcm5m3l1_ca_w_2_400_s_3_300 = 3.30e-05  mcm5m3l1_cc_w_2_400_s_3_300 = 9.10e-12  mcm5m3l1_cf_w_2_400_s_3_300 = 3.59e-11
+ mcm5m3l1_ca_w_2_400_s_9_000 = 3.30e-05  mcm5m3l1_cc_w_2_400_s_9_000 = 2.90e-13  mcm5m3l1_cf_w_2_400_s_9_000 = 4.40e-11
+ mcm5m3m1_ca_w_0_300_s_0_300 = 4.24e-05  mcm5m3m1_cc_w_0_300_s_0_300 = 8.40e-11  mcm5m3m1_cf_w_0_300_s_0_300 = 7.06e-12
+ mcm5m3m1_ca_w_0_300_s_0_360 = 4.24e-05  mcm5m3m1_cc_w_0_300_s_0_360 = 7.80e-11  mcm5m3m1_cf_w_0_300_s_0_360 = 8.25e-12
+ mcm5m3m1_ca_w_0_300_s_0_450 = 4.24e-05  mcm5m3m1_cc_w_0_300_s_0_450 = 6.98e-11  mcm5m3m1_cf_w_0_300_s_0_450 = 1.00e-11
+ mcm5m3m1_ca_w_0_300_s_0_600 = 4.24e-05  mcm5m3m1_cc_w_0_300_s_0_600 = 5.86e-11  mcm5m3m1_cf_w_0_300_s_0_600 = 1.29e-11
+ mcm5m3m1_ca_w_0_300_s_0_800 = 4.24e-05  mcm5m3m1_cc_w_0_300_s_0_800 = 4.71e-11  mcm5m3m1_cf_w_0_300_s_0_800 = 1.63e-11
+ mcm5m3m1_ca_w_0_300_s_1_000 = 4.24e-05  mcm5m3m1_cc_w_0_300_s_1_000 = 3.80e-11  mcm5m3m1_cf_w_0_300_s_1_000 = 1.95e-11
+ mcm5m3m1_ca_w_0_300_s_1_200 = 4.24e-05  mcm5m3m1_cc_w_0_300_s_1_200 = 3.12e-11  mcm5m3m1_cf_w_0_300_s_1_200 = 2.25e-11
+ mcm5m3m1_ca_w_0_300_s_2_100 = 4.24e-05  mcm5m3m1_cc_w_0_300_s_2_100 = 1.43e-11  mcm5m3m1_cf_w_0_300_s_2_100 = 3.26e-11
+ mcm5m3m1_ca_w_0_300_s_3_300 = 4.24e-05  mcm5m3m1_cc_w_0_300_s_3_300 = 5.57e-12  mcm5m3m1_cf_w_0_300_s_3_300 = 3.97e-11
+ mcm5m3m1_ca_w_0_300_s_9_000 = 4.24e-05  mcm5m3m1_cc_w_0_300_s_9_000 = 1.05e-13  mcm5m3m1_cf_w_0_300_s_9_000 = 4.49e-11
+ mcm5m3m1_ca_w_2_400_s_0_300 = 4.24e-05  mcm5m3m1_cc_w_2_400_s_0_300 = 9.41e-11  mcm5m3m1_cf_w_2_400_s_0_300 = 7.10e-12
+ mcm5m3m1_ca_w_2_400_s_0_360 = 4.24e-05  mcm5m3m1_cc_w_2_400_s_0_360 = 8.72e-11  mcm5m3m1_cf_w_2_400_s_0_360 = 8.28e-12
+ mcm5m3m1_ca_w_2_400_s_0_450 = 4.24e-05  mcm5m3m1_cc_w_2_400_s_0_450 = 7.77e-11  mcm5m3m1_cf_w_2_400_s_0_450 = 1.00e-11
+ mcm5m3m1_ca_w_2_400_s_0_600 = 4.24e-05  mcm5m3m1_cc_w_2_400_s_0_600 = 6.49e-11  mcm5m3m1_cf_w_2_400_s_0_600 = 1.28e-11
+ mcm5m3m1_ca_w_2_400_s_0_800 = 4.24e-05  mcm5m3m1_cc_w_2_400_s_0_800 = 5.20e-11  mcm5m3m1_cf_w_2_400_s_0_800 = 1.64e-11
+ mcm5m3m1_ca_w_2_400_s_1_000 = 4.24e-05  mcm5m3m1_cc_w_2_400_s_1_000 = 4.22e-11  mcm5m3m1_cf_w_2_400_s_1_000 = 1.97e-11
+ mcm5m3m1_ca_w_2_400_s_1_200 = 4.24e-05  mcm5m3m1_cc_w_2_400_s_1_200 = 3.48e-11  mcm5m3m1_cf_w_2_400_s_1_200 = 2.28e-11
+ mcm5m3m1_ca_w_2_400_s_2_100 = 4.24e-05  mcm5m3m1_cc_w_2_400_s_2_100 = 1.62e-11  mcm5m3m1_cf_w_2_400_s_2_100 = 3.35e-11
+ mcm5m3m1_ca_w_2_400_s_3_300 = 4.24e-05  mcm5m3m1_cc_w_2_400_s_3_300 = 6.39e-12  mcm5m3m1_cf_w_2_400_s_3_300 = 4.13e-11
+ mcm5m3m1_ca_w_2_400_s_9_000 = 4.24e-05  mcm5m3m1_cc_w_2_400_s_9_000 = 1.50e-13  mcm5m3m1_cf_w_2_400_s_9_000 = 4.71e-11
+ mcm5m3m2_ca_w_0_300_s_0_300 = 7.61e-05  mcm5m3m2_cc_w_0_300_s_0_300 = 7.79e-11  mcm5m3m2_cf_w_0_300_s_0_300 = 1.22e-11
+ mcm5m3m2_ca_w_0_300_s_0_360 = 7.61e-05  mcm5m3m2_cc_w_0_300_s_0_360 = 7.16e-11  mcm5m3m2_cf_w_0_300_s_0_360 = 1.41e-11
+ mcm5m3m2_ca_w_0_300_s_0_450 = 7.61e-05  mcm5m3m2_cc_w_0_300_s_0_450 = 6.30e-11  mcm5m3m2_cf_w_0_300_s_0_450 = 1.69e-11
+ mcm5m3m2_ca_w_0_300_s_0_600 = 7.61e-05  mcm5m3m2_cc_w_0_300_s_0_600 = 5.15e-11  mcm5m3m2_cf_w_0_300_s_0_600 = 2.13e-11
+ mcm5m3m2_ca_w_0_300_s_0_800 = 7.61e-05  mcm5m3m2_cc_w_0_300_s_0_800 = 3.97e-11  mcm5m3m2_cf_w_0_300_s_0_800 = 2.63e-11
+ mcm5m3m2_ca_w_0_300_s_1_000 = 7.61e-05  mcm5m3m2_cc_w_0_300_s_1_000 = 3.09e-11  mcm5m3m2_cf_w_0_300_s_1_000 = 3.08e-11
+ mcm5m3m2_ca_w_0_300_s_1_200 = 7.61e-05  mcm5m3m2_cc_w_0_300_s_1_200 = 2.43e-11  mcm5m3m2_cf_w_0_300_s_1_200 = 3.46e-11
+ mcm5m3m2_ca_w_0_300_s_2_100 = 7.61e-05  mcm5m3m2_cc_w_0_300_s_2_100 = 9.29e-12  mcm5m3m2_cf_w_0_300_s_2_100 = 4.57e-11
+ mcm5m3m2_ca_w_0_300_s_3_300 = 7.61e-05  mcm5m3m2_cc_w_0_300_s_3_300 = 2.92e-12  mcm5m3m2_cf_w_0_300_s_3_300 = 5.15e-11
+ mcm5m3m2_ca_w_0_300_s_9_000 = 7.61e-05  mcm5m3m2_cc_w_0_300_s_9_000 = 4.50e-14  mcm5m3m2_cf_w_0_300_s_9_000 = 5.43e-11
+ mcm5m3m2_ca_w_2_400_s_0_300 = 7.61e-05  mcm5m3m2_cc_w_2_400_s_0_300 = 8.49e-11  mcm5m3m2_cf_w_2_400_s_0_300 = 1.22e-11
+ mcm5m3m2_ca_w_2_400_s_0_360 = 7.61e-05  mcm5m3m2_cc_w_2_400_s_0_360 = 7.78e-11  mcm5m3m2_cf_w_2_400_s_0_360 = 1.42e-11
+ mcm5m3m2_ca_w_2_400_s_0_450 = 7.61e-05  mcm5m3m2_cc_w_2_400_s_0_450 = 6.88e-11  mcm5m3m2_cf_w_2_400_s_0_450 = 1.69e-11
+ mcm5m3m2_ca_w_2_400_s_0_600 = 7.61e-05  mcm5m3m2_cc_w_2_400_s_0_600 = 5.62e-11  mcm5m3m2_cf_w_2_400_s_0_600 = 2.13e-11
+ mcm5m3m2_ca_w_2_400_s_0_800 = 7.61e-05  mcm5m3m2_cc_w_2_400_s_0_800 = 4.35e-11  mcm5m3m2_cf_w_2_400_s_0_800 = 2.65e-11
+ mcm5m3m2_ca_w_2_400_s_1_000 = 7.61e-05  mcm5m3m2_cc_w_2_400_s_1_000 = 3.40e-11  mcm5m3m2_cf_w_2_400_s_1_000 = 3.10e-11
+ mcm5m3m2_ca_w_2_400_s_1_200 = 7.61e-05  mcm5m3m2_cc_w_2_400_s_1_200 = 2.70e-11  mcm5m3m2_cf_w_2_400_s_1_200 = 3.49e-11
+ mcm5m3m2_ca_w_2_400_s_2_100 = 7.61e-05  mcm5m3m2_cc_w_2_400_s_2_100 = 1.06e-11  mcm5m3m2_cf_w_2_400_s_2_100 = 4.66e-11
+ mcm5m3m2_ca_w_2_400_s_3_300 = 7.61e-05  mcm5m3m2_cc_w_2_400_s_3_300 = 3.41e-12  mcm5m3m2_cf_w_2_400_s_3_300 = 5.30e-11
+ mcm5m3m2_ca_w_2_400_s_9_000 = 7.61e-05  mcm5m3m2_cc_w_2_400_s_9_000 = 4.00e-14  mcm5m3m2_cf_w_2_400_s_9_000 = 5.63e-11
+ mcrdlm3f_ca_w_0_300_s_0_300 = 1.31e-05  mcrdlm3f_cc_w_0_300_s_0_300 = 9.14e-11  mcrdlm3f_cf_w_0_300_s_0_300 = 2.25e-12
+ mcrdlm3f_ca_w_0_300_s_0_360 = 1.31e-05  mcrdlm3f_cc_w_0_300_s_0_360 = 8.58e-11  mcrdlm3f_cf_w_0_300_s_0_360 = 2.64e-12
+ mcrdlm3f_ca_w_0_300_s_0_450 = 1.31e-05  mcrdlm3f_cc_w_0_300_s_0_450 = 7.81e-11  mcrdlm3f_cf_w_0_300_s_0_450 = 3.24e-12
+ mcrdlm3f_ca_w_0_300_s_0_600 = 1.31e-05  mcrdlm3f_cc_w_0_300_s_0_600 = 6.81e-11  mcrdlm3f_cf_w_0_300_s_0_600 = 4.22e-12
+ mcrdlm3f_ca_w_0_300_s_0_800 = 1.31e-05  mcrdlm3f_cc_w_0_300_s_0_800 = 5.81e-11  mcrdlm3f_cf_w_0_300_s_0_800 = 5.36e-12
+ mcrdlm3f_ca_w_0_300_s_1_000 = 1.31e-05  mcrdlm3f_cc_w_0_300_s_1_000 = 5.05e-11  mcrdlm3f_cf_w_0_300_s_1_000 = 6.55e-12
+ mcrdlm3f_ca_w_0_300_s_1_200 = 1.31e-05  mcrdlm3f_cc_w_0_300_s_1_200 = 4.46e-11  mcrdlm3f_cf_w_0_300_s_1_200 = 7.72e-12
+ mcrdlm3f_ca_w_0_300_s_2_100 = 1.31e-05  mcrdlm3f_cc_w_0_300_s_2_100 = 2.90e-11  mcrdlm3f_cf_w_0_300_s_2_100 = 1.27e-11
+ mcrdlm3f_ca_w_0_300_s_3_300 = 1.31e-05  mcrdlm3f_cc_w_0_300_s_3_300 = 1.93e-11  mcrdlm3f_cf_w_0_300_s_3_300 = 1.76e-11
+ mcrdlm3f_ca_w_0_300_s_9_000 = 1.31e-05  mcrdlm3f_cc_w_0_300_s_9_000 = 4.04e-12  mcrdlm3f_cf_w_0_300_s_9_000 = 2.89e-11
+ mcrdlm3f_ca_w_2_400_s_0_300 = 1.31e-05  mcrdlm3f_cc_w_2_400_s_0_300 = 1.15e-10  mcrdlm3f_cf_w_2_400_s_0_300 = 2.28e-12
+ mcrdlm3f_ca_w_2_400_s_0_360 = 1.31e-05  mcrdlm3f_cc_w_2_400_s_0_360 = 1.08e-10  mcrdlm3f_cf_w_2_400_s_0_360 = 2.67e-12
+ mcrdlm3f_ca_w_2_400_s_0_450 = 1.31e-05  mcrdlm3f_cc_w_2_400_s_0_450 = 9.90e-11  mcrdlm3f_cf_w_2_400_s_0_450 = 3.24e-12
+ mcrdlm3f_ca_w_2_400_s_0_600 = 1.31e-05  mcrdlm3f_cc_w_2_400_s_0_600 = 8.69e-11  mcrdlm3f_cf_w_2_400_s_0_600 = 4.18e-12
+ mcrdlm3f_ca_w_2_400_s_0_800 = 1.31e-05  mcrdlm3f_cc_w_2_400_s_0_800 = 7.44e-11  mcrdlm3f_cf_w_2_400_s_0_800 = 5.41e-12
+ mcrdlm3f_ca_w_2_400_s_1_000 = 1.31e-05  mcrdlm3f_cc_w_2_400_s_1_000 = 6.48e-11  mcrdlm3f_cf_w_2_400_s_1_000 = 6.62e-12
+ mcrdlm3f_ca_w_2_400_s_1_200 = 1.31e-05  mcrdlm3f_cc_w_2_400_s_1_200 = 5.74e-11  mcrdlm3f_cf_w_2_400_s_1_200 = 7.80e-12
+ mcrdlm3f_ca_w_2_400_s_2_100 = 1.31e-05  mcrdlm3f_cc_w_2_400_s_2_100 = 3.82e-11  mcrdlm3f_cf_w_2_400_s_2_100 = 1.27e-11
+ mcrdlm3f_ca_w_2_400_s_3_300 = 1.31e-05  mcrdlm3f_cc_w_2_400_s_3_300 = 2.54e-11  mcrdlm3f_cf_w_2_400_s_3_300 = 1.82e-11
+ mcrdlm3f_ca_w_2_400_s_9_000 = 1.31e-05  mcrdlm3f_cc_w_2_400_s_9_000 = 5.76e-12  mcrdlm3f_cf_w_2_400_s_9_000 = 3.20e-11
+ mcrdlm3d_ca_w_0_300_s_0_300 = 1.45e-05  mcrdlm3d_cc_w_0_300_s_0_300 = 9.12e-11  mcrdlm3d_cf_w_0_300_s_0_300 = 2.49e-12
+ mcrdlm3d_ca_w_0_300_s_0_360 = 1.45e-05  mcrdlm3d_cc_w_0_300_s_0_360 = 8.54e-11  mcrdlm3d_cf_w_0_300_s_0_360 = 2.92e-12
+ mcrdlm3d_ca_w_0_300_s_0_450 = 1.45e-05  mcrdlm3d_cc_w_0_300_s_0_450 = 7.77e-11  mcrdlm3d_cf_w_0_300_s_0_450 = 3.58e-12
+ mcrdlm3d_ca_w_0_300_s_0_600 = 1.45e-05  mcrdlm3d_cc_w_0_300_s_0_600 = 6.76e-11  mcrdlm3d_cf_w_0_300_s_0_600 = 4.66e-12
+ mcrdlm3d_ca_w_0_300_s_0_800 = 1.45e-05  mcrdlm3d_cc_w_0_300_s_0_800 = 5.75e-11  mcrdlm3d_cf_w_0_300_s_0_800 = 5.91e-12
+ mcrdlm3d_ca_w_0_300_s_1_000 = 1.45e-05  mcrdlm3d_cc_w_0_300_s_1_000 = 4.98e-11  mcrdlm3d_cf_w_0_300_s_1_000 = 7.22e-12
+ mcrdlm3d_ca_w_0_300_s_1_200 = 1.45e-05  mcrdlm3d_cc_w_0_300_s_1_200 = 4.39e-11  mcrdlm3d_cf_w_0_300_s_1_200 = 8.49e-12
+ mcrdlm3d_ca_w_0_300_s_2_100 = 1.45e-05  mcrdlm3d_cc_w_0_300_s_2_100 = 2.81e-11  mcrdlm3d_cf_w_0_300_s_2_100 = 1.39e-11
+ mcrdlm3d_ca_w_0_300_s_3_300 = 1.45e-05  mcrdlm3d_cc_w_0_300_s_3_300 = 1.83e-11  mcrdlm3d_cf_w_0_300_s_3_300 = 1.90e-11
+ mcrdlm3d_ca_w_0_300_s_9_000 = 1.45e-05  mcrdlm3d_cc_w_0_300_s_9_000 = 3.57e-12  mcrdlm3d_cf_w_0_300_s_9_000 = 3.03e-11
+ mcrdlm3d_ca_w_2_400_s_0_300 = 1.45e-05  mcrdlm3d_cc_w_2_400_s_0_300 = 1.14e-10  mcrdlm3d_cf_w_2_400_s_0_300 = 2.53e-12
+ mcrdlm3d_ca_w_2_400_s_0_360 = 1.45e-05  mcrdlm3d_cc_w_2_400_s_0_360 = 1.07e-10  mcrdlm3d_cf_w_2_400_s_0_360 = 2.95e-12
+ mcrdlm3d_ca_w_2_400_s_0_450 = 1.45e-05  mcrdlm3d_cc_w_2_400_s_0_450 = 9.78e-11  mcrdlm3d_cf_w_2_400_s_0_450 = 3.58e-12
+ mcrdlm3d_ca_w_2_400_s_0_600 = 1.45e-05  mcrdlm3d_cc_w_2_400_s_0_600 = 8.57e-11  mcrdlm3d_cf_w_2_400_s_0_600 = 4.62e-12
+ mcrdlm3d_ca_w_2_400_s_0_800 = 1.45e-05  mcrdlm3d_cc_w_2_400_s_0_800 = 7.32e-11  mcrdlm3d_cf_w_2_400_s_0_800 = 5.98e-12
+ mcrdlm3d_ca_w_2_400_s_1_000 = 1.45e-05  mcrdlm3d_cc_w_2_400_s_1_000 = 6.35e-11  mcrdlm3d_cf_w_2_400_s_1_000 = 7.30e-12
+ mcrdlm3d_ca_w_2_400_s_1_200 = 1.45e-05  mcrdlm3d_cc_w_2_400_s_1_200 = 5.61e-11  mcrdlm3d_cf_w_2_400_s_1_200 = 8.59e-12
+ mcrdlm3d_ca_w_2_400_s_2_100 = 1.45e-05  mcrdlm3d_cc_w_2_400_s_2_100 = 3.68e-11  mcrdlm3d_cf_w_2_400_s_2_100 = 1.39e-11
+ mcrdlm3d_ca_w_2_400_s_3_300 = 1.45e-05  mcrdlm3d_cc_w_2_400_s_3_300 = 2.41e-11  mcrdlm3d_cf_w_2_400_s_3_300 = 1.97e-11
+ mcrdlm3d_ca_w_2_400_s_9_000 = 1.45e-05  mcrdlm3d_cc_w_2_400_s_9_000 = 5.10e-12  mcrdlm3d_cf_w_2_400_s_9_000 = 3.36e-11
+ mcrdlm3p1_ca_w_0_300_s_0_300 = 1.55e-05  mcrdlm3p1_cc_w_0_300_s_0_300 = 9.09e-11  mcrdlm3p1_cf_w_0_300_s_0_300 = 2.66e-12
+ mcrdlm3p1_ca_w_0_300_s_0_360 = 1.55e-05  mcrdlm3p1_cc_w_0_300_s_0_360 = 8.49e-11  mcrdlm3p1_cf_w_0_300_s_0_360 = 3.12e-12
+ mcrdlm3p1_ca_w_0_300_s_0_450 = 1.55e-05  mcrdlm3p1_cc_w_0_300_s_0_450 = 7.74e-11  mcrdlm3p1_cf_w_0_300_s_0_450 = 3.82e-12
+ mcrdlm3p1_ca_w_0_300_s_0_600 = 1.55e-05  mcrdlm3p1_cc_w_0_300_s_0_600 = 6.72e-11  mcrdlm3p1_cf_w_0_300_s_0_600 = 4.96e-12
+ mcrdlm3p1_ca_w_0_300_s_0_800 = 1.55e-05  mcrdlm3p1_cc_w_0_300_s_0_800 = 5.71e-11  mcrdlm3p1_cf_w_0_300_s_0_800 = 6.28e-12
+ mcrdlm3p1_ca_w_0_300_s_1_000 = 1.55e-05  mcrdlm3p1_cc_w_0_300_s_1_000 = 4.94e-11  mcrdlm3p1_cf_w_0_300_s_1_000 = 7.68e-12
+ mcrdlm3p1_ca_w_0_300_s_1_200 = 1.55e-05  mcrdlm3p1_cc_w_0_300_s_1_200 = 4.34e-11  mcrdlm3p1_cf_w_0_300_s_1_200 = 9.02e-12
+ mcrdlm3p1_ca_w_0_300_s_2_100 = 1.55e-05  mcrdlm3p1_cc_w_0_300_s_2_100 = 2.75e-11  mcrdlm3p1_cf_w_0_300_s_2_100 = 1.47e-11
+ mcrdlm3p1_ca_w_0_300_s_3_300 = 1.55e-05  mcrdlm3p1_cc_w_0_300_s_3_300 = 1.77e-11  mcrdlm3p1_cf_w_0_300_s_3_300 = 2.00e-11
+ mcrdlm3p1_ca_w_0_300_s_9_000 = 1.55e-05  mcrdlm3p1_cc_w_0_300_s_9_000 = 3.30e-12  mcrdlm3p1_cf_w_0_300_s_9_000 = 3.12e-11
+ mcrdlm3p1_ca_w_2_400_s_0_300 = 1.55e-05  mcrdlm3p1_cc_w_2_400_s_0_300 = 1.13e-10  mcrdlm3p1_cf_w_2_400_s_0_300 = 2.72e-12
+ mcrdlm3p1_ca_w_2_400_s_0_360 = 1.55e-05  mcrdlm3p1_cc_w_2_400_s_0_360 = 1.06e-10  mcrdlm3p1_cf_w_2_400_s_0_360 = 3.17e-12
+ mcrdlm3p1_ca_w_2_400_s_0_450 = 1.55e-05  mcrdlm3p1_cc_w_2_400_s_0_450 = 9.71e-11  mcrdlm3p1_cf_w_2_400_s_0_450 = 3.84e-12
+ mcrdlm3p1_ca_w_2_400_s_0_600 = 1.55e-05  mcrdlm3p1_cc_w_2_400_s_0_600 = 8.49e-11  mcrdlm3p1_cf_w_2_400_s_0_600 = 4.95e-12
+ mcrdlm3p1_ca_w_2_400_s_0_800 = 1.55e-05  mcrdlm3p1_cc_w_2_400_s_0_800 = 7.24e-11  mcrdlm3p1_cf_w_2_400_s_0_800 = 6.38e-12
+ mcrdlm3p1_ca_w_2_400_s_1_000 = 1.55e-05  mcrdlm3p1_cc_w_2_400_s_1_000 = 6.26e-11  mcrdlm3p1_cf_w_2_400_s_1_000 = 7.79e-12
+ mcrdlm3p1_ca_w_2_400_s_1_200 = 1.55e-05  mcrdlm3p1_cc_w_2_400_s_1_200 = 5.54e-11  mcrdlm3p1_cf_w_2_400_s_1_200 = 9.15e-12
+ mcrdlm3p1_ca_w_2_400_s_2_100 = 1.55e-05  mcrdlm3p1_cc_w_2_400_s_2_100 = 3.60e-11  mcrdlm3p1_cf_w_2_400_s_2_100 = 1.47e-11
+ mcrdlm3p1_ca_w_2_400_s_3_300 = 1.55e-05  mcrdlm3p1_cc_w_2_400_s_3_300 = 2.34e-11  mcrdlm3p1_cf_w_2_400_s_3_300 = 2.08e-11
+ mcrdlm3p1_ca_w_2_400_s_9_000 = 1.55e-05  mcrdlm3p1_cc_w_2_400_s_9_000 = 4.77e-12  mcrdlm3p1_cf_w_2_400_s_9_000 = 3.46e-11
+ mcrdlm3l1_ca_w_0_300_s_0_300 = 1.92e-05  mcrdlm3l1_cc_w_0_300_s_0_300 = 9.00e-11  mcrdlm3l1_cf_w_0_300_s_0_300 = 3.27e-12
+ mcrdlm3l1_ca_w_0_300_s_0_360 = 1.92e-05  mcrdlm3l1_cc_w_0_300_s_0_360 = 8.40e-11  mcrdlm3l1_cf_w_0_300_s_0_360 = 3.82e-12
+ mcrdlm3l1_ca_w_0_300_s_0_450 = 1.92e-05  mcrdlm3l1_cc_w_0_300_s_0_450 = 7.67e-11  mcrdlm3l1_cf_w_0_300_s_0_450 = 4.67e-12
+ mcrdlm3l1_ca_w_0_300_s_0_600 = 1.92e-05  mcrdlm3l1_cc_w_0_300_s_0_600 = 6.60e-11  mcrdlm3l1_cf_w_0_300_s_0_600 = 6.04e-12
+ mcrdlm3l1_ca_w_0_300_s_0_800 = 1.92e-05  mcrdlm3l1_cc_w_0_300_s_0_800 = 5.56e-11  mcrdlm3l1_cf_w_0_300_s_0_800 = 7.68e-12
+ mcrdlm3l1_ca_w_0_300_s_1_000 = 1.92e-05  mcrdlm3l1_cc_w_0_300_s_1_000 = 4.78e-11  mcrdlm3l1_cf_w_0_300_s_1_000 = 9.33e-12
+ mcrdlm3l1_ca_w_0_300_s_1_200 = 1.92e-05  mcrdlm3l1_cc_w_0_300_s_1_200 = 4.17e-11  mcrdlm3l1_cf_w_0_300_s_1_200 = 1.09e-11
+ mcrdlm3l1_ca_w_0_300_s_2_100 = 1.92e-05  mcrdlm3l1_cc_w_0_300_s_2_100 = 2.56e-11  mcrdlm3l1_cf_w_0_300_s_2_100 = 1.74e-11
+ mcrdlm3l1_ca_w_0_300_s_3_300 = 1.92e-05  mcrdlm3l1_cc_w_0_300_s_3_300 = 1.58e-11  mcrdlm3l1_cf_w_0_300_s_3_300 = 2.32e-11
+ mcrdlm3l1_ca_w_0_300_s_9_000 = 1.92e-05  mcrdlm3l1_cc_w_0_300_s_9_000 = 2.58e-12  mcrdlm3l1_cf_w_0_300_s_9_000 = 3.41e-11
+ mcrdlm3l1_ca_w_2_400_s_0_300 = 1.92e-05  mcrdlm3l1_cc_w_2_400_s_0_300 = 1.11e-10  mcrdlm3l1_cf_w_2_400_s_0_300 = 3.31e-12
+ mcrdlm3l1_ca_w_2_400_s_0_360 = 1.92e-05  mcrdlm3l1_cc_w_2_400_s_0_360 = 1.04e-10  mcrdlm3l1_cf_w_2_400_s_0_360 = 3.85e-12
+ mcrdlm3l1_ca_w_2_400_s_0_450 = 1.92e-05  mcrdlm3l1_cc_w_2_400_s_0_450 = 9.45e-11  mcrdlm3l1_cf_w_2_400_s_0_450 = 4.67e-12
+ mcrdlm3l1_ca_w_2_400_s_0_600 = 1.92e-05  mcrdlm3l1_cc_w_2_400_s_0_600 = 8.23e-11  mcrdlm3l1_cf_w_2_400_s_0_600 = 6.02e-12
+ mcrdlm3l1_ca_w_2_400_s_0_800 = 1.92e-05  mcrdlm3l1_cc_w_2_400_s_0_800 = 6.97e-11  mcrdlm3l1_cf_w_2_400_s_0_800 = 7.75e-12
+ mcrdlm3l1_ca_w_2_400_s_1_000 = 1.92e-05  mcrdlm3l1_cc_w_2_400_s_1_000 = 6.00e-11  mcrdlm3l1_cf_w_2_400_s_1_000 = 9.44e-12
+ mcrdlm3l1_ca_w_2_400_s_1_200 = 1.92e-05  mcrdlm3l1_cc_w_2_400_s_1_200 = 5.27e-11  mcrdlm3l1_cf_w_2_400_s_1_200 = 1.10e-11
+ mcrdlm3l1_ca_w_2_400_s_2_100 = 1.92e-05  mcrdlm3l1_cc_w_2_400_s_2_100 = 3.35e-11  mcrdlm3l1_cf_w_2_400_s_2_100 = 1.75e-11
+ mcrdlm3l1_ca_w_2_400_s_3_300 = 1.92e-05  mcrdlm3l1_cc_w_2_400_s_3_300 = 2.11e-11  mcrdlm3l1_cf_w_2_400_s_3_300 = 2.42e-11
+ mcrdlm3l1_ca_w_2_400_s_9_000 = 1.92e-05  mcrdlm3l1_cc_w_2_400_s_9_000 = 3.85e-12  mcrdlm3l1_cf_w_2_400_s_9_000 = 3.78e-11
+ mcrdlm3m1_ca_w_0_300_s_0_300 = 2.87e-05  mcrdlm3m1_cc_w_0_300_s_0_300 = 8.76e-11  mcrdlm3m1_cf_w_0_300_s_0_300 = 4.80e-12
+ mcrdlm3m1_ca_w_0_300_s_0_360 = 2.87e-05  mcrdlm3m1_cc_w_0_300_s_0_360 = 8.17e-11  mcrdlm3m1_cf_w_0_300_s_0_360 = 5.60e-12
+ mcrdlm3m1_ca_w_0_300_s_0_450 = 2.87e-05  mcrdlm3m1_cc_w_0_300_s_0_450 = 7.40e-11  mcrdlm3m1_cf_w_0_300_s_0_450 = 6.80e-12
+ mcrdlm3m1_ca_w_0_300_s_0_600 = 2.87e-05  mcrdlm3m1_cc_w_0_300_s_0_600 = 6.32e-11  mcrdlm3m1_cf_w_0_300_s_0_600 = 8.73e-12
+ mcrdlm3m1_ca_w_0_300_s_0_800 = 2.87e-05  mcrdlm3m1_cc_w_0_300_s_0_800 = 5.24e-11  mcrdlm3m1_cf_w_0_300_s_0_800 = 1.11e-11
+ mcrdlm3m1_ca_w_0_300_s_1_000 = 2.87e-05  mcrdlm3m1_cc_w_0_300_s_1_000 = 4.44e-11  mcrdlm3m1_cf_w_0_300_s_1_000 = 1.33e-11
+ mcrdlm3m1_ca_w_0_300_s_1_200 = 2.87e-05  mcrdlm3m1_cc_w_0_300_s_1_200 = 3.81e-11  mcrdlm3m1_cf_w_0_300_s_1_200 = 1.54e-11
+ mcrdlm3m1_ca_w_0_300_s_2_100 = 2.87e-05  mcrdlm3m1_cc_w_0_300_s_2_100 = 2.18e-11  mcrdlm3m1_cf_w_0_300_s_2_100 = 2.36e-11
+ mcrdlm3m1_ca_w_0_300_s_3_300 = 2.87e-05  mcrdlm3m1_cc_w_0_300_s_3_300 = 1.25e-11  mcrdlm3m1_cf_w_0_300_s_3_300 = 3.00e-11
+ mcrdlm3m1_ca_w_0_300_s_9_000 = 2.87e-05  mcrdlm3m1_cc_w_0_300_s_9_000 = 1.69e-12  mcrdlm3m1_cf_w_0_300_s_9_000 = 3.95e-11
+ mcrdlm3m1_ca_w_2_400_s_0_300 = 2.87e-05  mcrdlm3m1_cc_w_2_400_s_0_300 = 1.06e-10  mcrdlm3m1_cf_w_2_400_s_0_300 = 4.82e-12
+ mcrdlm3m1_ca_w_2_400_s_0_360 = 2.87e-05  mcrdlm3m1_cc_w_2_400_s_0_360 = 9.87e-11  mcrdlm3m1_cf_w_2_400_s_0_360 = 5.62e-12
+ mcrdlm3m1_ca_w_2_400_s_0_450 = 2.87e-05  mcrdlm3m1_cc_w_2_400_s_0_450 = 8.97e-11  mcrdlm3m1_cf_w_2_400_s_0_450 = 6.80e-12
+ mcrdlm3m1_ca_w_2_400_s_0_600 = 2.87e-05  mcrdlm3m1_cc_w_2_400_s_0_600 = 7.74e-11  mcrdlm3m1_cf_w_2_400_s_0_600 = 8.70e-12
+ mcrdlm3m1_ca_w_2_400_s_0_800 = 2.87e-05  mcrdlm3m1_cc_w_2_400_s_0_800 = 6.49e-11  mcrdlm3m1_cf_w_2_400_s_0_800 = 1.11e-11
+ mcrdlm3m1_ca_w_2_400_s_1_000 = 2.87e-05  mcrdlm3m1_cc_w_2_400_s_1_000 = 5.53e-11  mcrdlm3m1_cf_w_2_400_s_1_000 = 1.34e-11
+ mcrdlm3m1_ca_w_2_400_s_1_200 = 2.87e-05  mcrdlm3m1_cc_w_2_400_s_1_200 = 4.79e-11  mcrdlm3m1_cf_w_2_400_s_1_200 = 1.56e-11
+ mcrdlm3m1_ca_w_2_400_s_2_100 = 2.87e-05  mcrdlm3m1_cc_w_2_400_s_2_100 = 2.90e-11  mcrdlm3m1_cf_w_2_400_s_2_100 = 2.37e-11
+ mcrdlm3m1_ca_w_2_400_s_3_300 = 2.87e-05  mcrdlm3m1_cc_w_2_400_s_3_300 = 1.74e-11  mcrdlm3m1_cf_w_2_400_s_3_300 = 3.13e-11
+ mcrdlm3m1_ca_w_2_400_s_9_000 = 2.87e-05  mcrdlm3m1_cc_w_2_400_s_9_000 = 2.68e-12  mcrdlm3m1_cf_w_2_400_s_9_000 = 4.37e-11
+ mcrdlm3m2_ca_w_0_300_s_0_300 = 6.23e-05  mcrdlm3m2_cc_w_0_300_s_0_300 = 8.15e-11  mcrdlm3m2_cf_w_0_300_s_0_300 = 9.93e-12
+ mcrdlm3m2_ca_w_0_300_s_0_360 = 6.23e-05  mcrdlm3m2_cc_w_0_300_s_0_360 = 7.51e-11  mcrdlm3m2_cf_w_0_300_s_0_360 = 1.15e-11
+ mcrdlm3m2_ca_w_0_300_s_0_450 = 6.23e-05  mcrdlm3m2_cc_w_0_300_s_0_450 = 6.73e-11  mcrdlm3m2_cf_w_0_300_s_0_450 = 1.37e-11
+ mcrdlm3m2_ca_w_0_300_s_0_600 = 6.23e-05  mcrdlm3m2_cc_w_0_300_s_0_600 = 5.62e-11  mcrdlm3m2_cf_w_0_300_s_0_600 = 1.72e-11
+ mcrdlm3m2_ca_w_0_300_s_0_800 = 6.23e-05  mcrdlm3m2_cc_w_0_300_s_0_800 = 4.53e-11  mcrdlm3m2_cf_w_0_300_s_0_800 = 2.12e-11
+ mcrdlm3m2_ca_w_0_300_s_1_000 = 6.23e-05  mcrdlm3m2_cc_w_0_300_s_1_000 = 3.70e-11  mcrdlm3m2_cf_w_0_300_s_1_000 = 2.48e-11
+ mcrdlm3m2_ca_w_0_300_s_1_200 = 6.23e-05  mcrdlm3m2_cc_w_0_300_s_1_200 = 3.10e-11  mcrdlm3m2_cf_w_0_300_s_1_200 = 2.79e-11
+ mcrdlm3m2_ca_w_0_300_s_2_100 = 6.23e-05  mcrdlm3m2_cc_w_0_300_s_2_100 = 1.55e-11  mcrdlm3m2_cf_w_0_300_s_2_100 = 3.82e-11
+ mcrdlm3m2_ca_w_0_300_s_3_300 = 6.23e-05  mcrdlm3m2_cc_w_0_300_s_3_300 = 8.00e-12  mcrdlm3m2_cf_w_0_300_s_3_300 = 4.46e-11
+ mcrdlm3m2_ca_w_0_300_s_9_000 = 6.23e-05  mcrdlm3m2_cc_w_0_300_s_9_000 = 8.83e-13  mcrdlm3m2_cf_w_0_300_s_9_000 = 5.13e-11
+ mcrdlm3m2_ca_w_2_400_s_0_300 = 6.23e-05  mcrdlm3m2_cc_w_2_400_s_0_300 = 9.66e-11  mcrdlm3m2_cf_w_2_400_s_0_300 = 9.96e-12
+ mcrdlm3m2_ca_w_2_400_s_0_360 = 6.23e-05  mcrdlm3m2_cc_w_2_400_s_0_360 = 8.97e-11  mcrdlm3m2_cf_w_2_400_s_0_360 = 1.15e-11
+ mcrdlm3m2_ca_w_2_400_s_0_450 = 6.23e-05  mcrdlm3m2_cc_w_2_400_s_0_450 = 8.08e-11  mcrdlm3m2_cf_w_2_400_s_0_450 = 1.37e-11
+ mcrdlm3m2_ca_w_2_400_s_0_600 = 6.23e-05  mcrdlm3m2_cc_w_2_400_s_0_600 = 6.87e-11  mcrdlm3m2_cf_w_2_400_s_0_600 = 1.72e-11
+ mcrdlm3m2_ca_w_2_400_s_0_800 = 6.23e-05  mcrdlm3m2_cc_w_2_400_s_0_800 = 5.62e-11  mcrdlm3m2_cf_w_2_400_s_0_800 = 2.13e-11
+ mcrdlm3m2_ca_w_2_400_s_1_000 = 6.23e-05  mcrdlm3m2_cc_w_2_400_s_1_000 = 4.70e-11  mcrdlm3m2_cf_w_2_400_s_1_000 = 2.49e-11
+ mcrdlm3m2_ca_w_2_400_s_1_200 = 6.23e-05  mcrdlm3m2_cc_w_2_400_s_1_200 = 4.00e-11  mcrdlm3m2_cf_w_2_400_s_1_200 = 2.82e-11
+ mcrdlm3m2_ca_w_2_400_s_2_100 = 6.23e-05  mcrdlm3m2_cc_w_2_400_s_2_100 = 2.25e-11  mcrdlm3m2_cf_w_2_400_s_2_100 = 3.86e-11
+ mcrdlm3m2_ca_w_2_400_s_3_300 = 6.23e-05  mcrdlm3m2_cc_w_2_400_s_3_300 = 1.25e-11  mcrdlm3m2_cf_w_2_400_s_3_300 = 4.65e-11
+ mcrdlm3m2_ca_w_2_400_s_9_000 = 6.23e-05  mcrdlm3m2_cc_w_2_400_s_9_000 = 1.67e-12  mcrdlm3m2_cf_w_2_400_s_9_000 = 5.65e-11
+ mcm5m4f_ca_w_0_300_s_0_300 = 5.59e-05  mcm5m4f_cc_w_0_300_s_0_300 = 8.25e-11  mcm5m4f_cf_w_0_300_s_0_300 = 8.68e-12
+ mcm5m4f_ca_w_0_300_s_0_360 = 5.59e-05  mcm5m4f_cc_w_0_300_s_0_360 = 7.61e-11  mcm5m4f_cf_w_0_300_s_0_360 = 1.01e-11
+ mcm5m4f_ca_w_0_300_s_0_450 = 5.59e-05  mcm5m4f_cc_w_0_300_s_0_450 = 6.78e-11  mcm5m4f_cf_w_0_300_s_0_450 = 1.22e-11
+ mcm5m4f_ca_w_0_300_s_0_600 = 5.59e-05  mcm5m4f_cc_w_0_300_s_0_600 = 5.67e-11  mcm5m4f_cf_w_0_300_s_0_600 = 1.55e-11
+ mcm5m4f_ca_w_0_300_s_0_800 = 5.59e-05  mcm5m4f_cc_w_0_300_s_0_800 = 4.54e-11  mcm5m4f_cf_w_0_300_s_0_800 = 1.94e-11
+ mcm5m4f_ca_w_0_300_s_1_000 = 5.59e-05  mcm5m4f_cc_w_0_300_s_1_000 = 3.70e-11  mcm5m4f_cf_w_0_300_s_1_000 = 2.29e-11
+ mcm5m4f_ca_w_0_300_s_1_200 = 5.59e-05  mcm5m4f_cc_w_0_300_s_1_200 = 3.05e-11  mcm5m4f_cf_w_0_300_s_1_200 = 2.60e-11
+ mcm5m4f_ca_w_0_300_s_2_100 = 5.59e-05  mcm5m4f_cc_w_0_300_s_2_100 = 1.45e-11  mcm5m4f_cf_w_0_300_s_2_100 = 3.63e-11
+ mcm5m4f_ca_w_0_300_s_3_300 = 5.59e-05  mcm5m4f_cc_w_0_300_s_3_300 = 6.47e-12  mcm5m4f_cf_w_0_300_s_3_300 = 4.30e-11
+ mcm5m4f_ca_w_0_300_s_9_000 = 5.59e-05  mcm5m4f_cc_w_0_300_s_9_000 = 3.00e-13  mcm5m4f_cf_w_0_300_s_9_000 = 4.88e-11
+ mcm5m4f_ca_w_2_400_s_0_300 = 5.59e-05  mcm5m4f_cc_w_2_400_s_0_300 = 9.44e-11  mcm5m4f_cf_w_2_400_s_0_300 = 8.76e-12
+ mcm5m4f_ca_w_2_400_s_0_360 = 5.59e-05  mcm5m4f_cc_w_2_400_s_0_360 = 8.75e-11  mcm5m4f_cf_w_2_400_s_0_360 = 1.02e-11
+ mcm5m4f_ca_w_2_400_s_0_450 = 5.59e-05  mcm5m4f_cc_w_2_400_s_0_450 = 7.86e-11  mcm5m4f_cf_w_2_400_s_0_450 = 1.23e-11
+ mcm5m4f_ca_w_2_400_s_0_600 = 5.59e-05  mcm5m4f_cc_w_2_400_s_0_600 = 6.59e-11  mcm5m4f_cf_w_2_400_s_0_600 = 1.55e-11
+ mcm5m4f_ca_w_2_400_s_0_800 = 5.59e-05  mcm5m4f_cc_w_2_400_s_0_800 = 5.32e-11  mcm5m4f_cf_w_2_400_s_0_800 = 1.96e-11
+ mcm5m4f_ca_w_2_400_s_1_000 = 5.59e-05  mcm5m4f_cc_w_2_400_s_1_000 = 4.36e-11  mcm5m4f_cf_w_2_400_s_1_000 = 2.32e-11
+ mcm5m4f_ca_w_2_400_s_1_200 = 5.59e-05  mcm5m4f_cc_w_2_400_s_1_200 = 3.64e-11  mcm5m4f_cf_w_2_400_s_1_200 = 2.64e-11
+ mcm5m4f_ca_w_2_400_s_2_100 = 5.59e-05  mcm5m4f_cc_w_2_400_s_2_100 = 1.85e-11  mcm5m4f_cf_w_2_400_s_2_100 = 3.71e-11
+ mcm5m4f_ca_w_2_400_s_3_300 = 5.59e-05  mcm5m4f_cc_w_2_400_s_3_300 = 8.71e-12  mcm5m4f_cf_w_2_400_s_3_300 = 4.48e-11
+ mcm5m4f_ca_w_2_400_s_9_000 = 5.59e-05  mcm5m4f_cc_w_2_400_s_9_000 = 4.30e-13  mcm5m4f_cf_w_2_400_s_9_000 = 5.26e-11
+ mcm5m4d_ca_w_0_300_s_0_300 = 5.66e-05  mcm5m4d_cc_w_0_300_s_0_300 = 8.23e-11  mcm5m4d_cf_w_0_300_s_0_300 = 8.80e-12
+ mcm5m4d_ca_w_0_300_s_0_360 = 5.66e-05  mcm5m4d_cc_w_0_300_s_0_360 = 7.59e-11  mcm5m4d_cf_w_0_300_s_0_360 = 1.02e-11
+ mcm5m4d_ca_w_0_300_s_0_450 = 5.66e-05  mcm5m4d_cc_w_0_300_s_0_450 = 6.76e-11  mcm5m4d_cf_w_0_300_s_0_450 = 1.24e-11
+ mcm5m4d_ca_w_0_300_s_0_600 = 5.66e-05  mcm5m4d_cc_w_0_300_s_0_600 = 5.65e-11  mcm5m4d_cf_w_0_300_s_0_600 = 1.57e-11
+ mcm5m4d_ca_w_0_300_s_0_800 = 5.66e-05  mcm5m4d_cc_w_0_300_s_0_800 = 4.51e-11  mcm5m4d_cf_w_0_300_s_0_800 = 1.96e-11
+ mcm5m4d_ca_w_0_300_s_1_000 = 5.66e-05  mcm5m4d_cc_w_0_300_s_1_000 = 3.66e-11  mcm5m4d_cf_w_0_300_s_1_000 = 2.32e-11
+ mcm5m4d_ca_w_0_300_s_1_200 = 5.66e-05  mcm5m4d_cc_w_0_300_s_1_200 = 3.01e-11  mcm5m4d_cf_w_0_300_s_1_200 = 2.64e-11
+ mcm5m4d_ca_w_0_300_s_2_100 = 5.66e-05  mcm5m4d_cc_w_0_300_s_2_100 = 1.41e-11  mcm5m4d_cf_w_0_300_s_2_100 = 3.67e-11
+ mcm5m4d_ca_w_0_300_s_3_300 = 5.66e-05  mcm5m4d_cc_w_0_300_s_3_300 = 6.18e-12  mcm5m4d_cf_w_0_300_s_3_300 = 4.34e-11
+ mcm5m4d_ca_w_0_300_s_9_000 = 5.66e-05  mcm5m4d_cc_w_0_300_s_9_000 = 2.40e-13  mcm5m4d_cf_w_0_300_s_9_000 = 4.89e-11
+ mcm5m4d_ca_w_2_400_s_0_300 = 5.66e-05  mcm5m4d_cc_w_2_400_s_0_300 = 9.37e-11  mcm5m4d_cf_w_2_400_s_0_300 = 8.88e-12
+ mcm5m4d_ca_w_2_400_s_0_360 = 5.66e-05  mcm5m4d_cc_w_2_400_s_0_360 = 8.68e-11  mcm5m4d_cf_w_2_400_s_0_360 = 1.03e-11
+ mcm5m4d_ca_w_2_400_s_0_450 = 5.66e-05  mcm5m4d_cc_w_2_400_s_0_450 = 7.79e-11  mcm5m4d_cf_w_2_400_s_0_450 = 1.24e-11
+ mcm5m4d_ca_w_2_400_s_0_600 = 5.66e-05  mcm5m4d_cc_w_2_400_s_0_600 = 6.52e-11  mcm5m4d_cf_w_2_400_s_0_600 = 1.58e-11
+ mcm5m4d_ca_w_2_400_s_0_800 = 5.66e-05  mcm5m4d_cc_w_2_400_s_0_800 = 5.25e-11  mcm5m4d_cf_w_2_400_s_0_800 = 1.98e-11
+ mcm5m4d_ca_w_2_400_s_1_000 = 5.66e-05  mcm5m4d_cc_w_2_400_s_1_000 = 4.29e-11  mcm5m4d_cf_w_2_400_s_1_000 = 2.35e-11
+ mcm5m4d_ca_w_2_400_s_1_200 = 5.66e-05  mcm5m4d_cc_w_2_400_s_1_200 = 3.56e-11  mcm5m4d_cf_w_2_400_s_1_200 = 2.68e-11
+ mcm5m4d_ca_w_2_400_s_2_100 = 5.66e-05  mcm5m4d_cc_w_2_400_s_2_100 = 1.78e-11  mcm5m4d_cf_w_2_400_s_2_100 = 3.75e-11
+ mcm5m4d_ca_w_2_400_s_3_300 = 5.66e-05  mcm5m4d_cc_w_2_400_s_3_300 = 8.15e-12  mcm5m4d_cf_w_2_400_s_3_300 = 4.52e-11
+ mcm5m4d_ca_w_2_400_s_9_000 = 5.66e-05  mcm5m4d_cc_w_2_400_s_9_000 = 3.95e-13  mcm5m4d_cf_w_2_400_s_9_000 = 5.25e-11
+ mcm5m4p1_ca_w_0_300_s_0_300 = 5.71e-05  mcm5m4p1_cc_w_0_300_s_0_300 = 8.20e-11  mcm5m4p1_cf_w_0_300_s_0_300 = 8.87e-12
+ mcm5m4p1_ca_w_0_300_s_0_360 = 5.71e-05  mcm5m4p1_cc_w_0_300_s_0_360 = 7.58e-11  mcm5m4p1_cf_w_0_300_s_0_360 = 1.03e-11
+ mcm5m4p1_ca_w_0_300_s_0_450 = 5.71e-05  mcm5m4p1_cc_w_0_300_s_0_450 = 6.75e-11  mcm5m4p1_cf_w_0_300_s_0_450 = 1.25e-11
+ mcm5m4p1_ca_w_0_300_s_0_600 = 5.71e-05  mcm5m4p1_cc_w_0_300_s_0_600 = 5.63e-11  mcm5m4p1_cf_w_0_300_s_0_600 = 1.59e-11
+ mcm5m4p1_ca_w_0_300_s_0_800 = 5.71e-05  mcm5m4p1_cc_w_0_300_s_0_800 = 4.49e-11  mcm5m4p1_cf_w_0_300_s_0_800 = 1.98e-11
+ mcm5m4p1_ca_w_0_300_s_1_000 = 5.71e-05  mcm5m4p1_cc_w_0_300_s_1_000 = 3.64e-11  mcm5m4p1_cf_w_0_300_s_1_000 = 2.34e-11
+ mcm5m4p1_ca_w_0_300_s_1_200 = 5.71e-05  mcm5m4p1_cc_w_0_300_s_1_200 = 2.99e-11  mcm5m4p1_cf_w_0_300_s_1_200 = 2.66e-11
+ mcm5m4p1_ca_w_0_300_s_2_100 = 5.71e-05  mcm5m4p1_cc_w_0_300_s_2_100 = 1.39e-11  mcm5m4p1_cf_w_0_300_s_2_100 = 3.70e-11
+ mcm5m4p1_ca_w_0_300_s_3_300 = 5.71e-05  mcm5m4p1_cc_w_0_300_s_3_300 = 5.96e-12  mcm5m4p1_cf_w_0_300_s_3_300 = 4.36e-11
+ mcm5m4p1_ca_w_0_300_s_9_000 = 5.71e-05  mcm5m4p1_cc_w_0_300_s_9_000 = 2.45e-13  mcm5m4p1_cf_w_0_300_s_9_000 = 4.91e-11
+ mcm5m4p1_ca_w_2_400_s_0_300 = 5.71e-05  mcm5m4p1_cc_w_2_400_s_0_300 = 9.32e-11  mcm5m4p1_cf_w_2_400_s_0_300 = 8.96e-12
+ mcm5m4p1_ca_w_2_400_s_0_360 = 5.71e-05  mcm5m4p1_cc_w_2_400_s_0_360 = 8.65e-11  mcm5m4p1_cf_w_2_400_s_0_360 = 1.04e-11
+ mcm5m4p1_ca_w_2_400_s_0_450 = 5.71e-05  mcm5m4p1_cc_w_2_400_s_0_450 = 7.73e-11  mcm5m4p1_cf_w_2_400_s_0_450 = 1.25e-11
+ mcm5m4p1_ca_w_2_400_s_0_600 = 5.71e-05  mcm5m4p1_cc_w_2_400_s_0_600 = 6.47e-11  mcm5m4p1_cf_w_2_400_s_0_600 = 1.59e-11
+ mcm5m4p1_ca_w_2_400_s_0_800 = 5.71e-05  mcm5m4p1_cc_w_2_400_s_0_800 = 5.20e-11  mcm5m4p1_cf_w_2_400_s_0_800 = 2.00e-11
+ mcm5m4p1_ca_w_2_400_s_1_000 = 5.71e-05  mcm5m4p1_cc_w_2_400_s_1_000 = 4.24e-11  mcm5m4p1_cf_w_2_400_s_1_000 = 2.37e-11
+ mcm5m4p1_ca_w_2_400_s_1_200 = 5.71e-05  mcm5m4p1_cc_w_2_400_s_1_200 = 3.52e-11  mcm5m4p1_cf_w_2_400_s_1_200 = 2.70e-11
+ mcm5m4p1_ca_w_2_400_s_2_100 = 5.71e-05  mcm5m4p1_cc_w_2_400_s_2_100 = 1.73e-11  mcm5m4p1_cf_w_2_400_s_2_100 = 3.78e-11
+ mcm5m4p1_ca_w_2_400_s_3_300 = 5.71e-05  mcm5m4p1_cc_w_2_400_s_3_300 = 7.77e-12  mcm5m4p1_cf_w_2_400_s_3_300 = 4.55e-11
+ mcm5m4p1_ca_w_2_400_s_9_000 = 5.71e-05  mcm5m4p1_cc_w_2_400_s_9_000 = 3.60e-13  mcm5m4p1_cf_w_2_400_s_9_000 = 5.25e-11
+ mcm5m4l1_ca_w_0_300_s_0_300 = 5.86e-05  mcm5m4l1_cc_w_0_300_s_0_300 = 8.16e-11  mcm5m4l1_cf_w_0_300_s_0_300 = 9.12e-12
+ mcm5m4l1_ca_w_0_300_s_0_360 = 5.86e-05  mcm5m4l1_cc_w_0_300_s_0_360 = 7.53e-11  mcm5m4l1_cf_w_0_300_s_0_360 = 1.06e-11
+ mcm5m4l1_ca_w_0_300_s_0_450 = 5.86e-05  mcm5m4l1_cc_w_0_300_s_0_450 = 6.72e-11  mcm5m4l1_cf_w_0_300_s_0_450 = 1.28e-11
+ mcm5m4l1_ca_w_0_300_s_0_600 = 5.86e-05  mcm5m4l1_cc_w_0_300_s_0_600 = 5.58e-11  mcm5m4l1_cf_w_0_300_s_0_600 = 1.63e-11
+ mcm5m4l1_ca_w_0_300_s_0_800 = 5.86e-05  mcm5m4l1_cc_w_0_300_s_0_800 = 4.43e-11  mcm5m4l1_cf_w_0_300_s_0_800 = 2.04e-11
+ mcm5m4l1_ca_w_0_300_s_1_000 = 5.86e-05  mcm5m4l1_cc_w_0_300_s_1_000 = 3.57e-11  mcm5m4l1_cf_w_0_300_s_1_000 = 2.41e-11
+ mcm5m4l1_ca_w_0_300_s_1_200 = 5.86e-05  mcm5m4l1_cc_w_0_300_s_1_200 = 2.92e-11  mcm5m4l1_cf_w_0_300_s_1_200 = 2.74e-11
+ mcm5m4l1_ca_w_0_300_s_2_100 = 5.86e-05  mcm5m4l1_cc_w_0_300_s_2_100 = 1.32e-11  mcm5m4l1_cf_w_0_300_s_2_100 = 3.78e-11
+ mcm5m4l1_ca_w_0_300_s_3_300 = 5.86e-05  mcm5m4l1_cc_w_0_300_s_3_300 = 5.35e-12  mcm5m4l1_cf_w_0_300_s_3_300 = 4.44e-11
+ mcm5m4l1_ca_w_0_300_s_9_000 = 5.86e-05  mcm5m4l1_cc_w_0_300_s_9_000 = 1.80e-13  mcm5m4l1_cf_w_0_300_s_9_000 = 4.94e-11
+ mcm5m4l1_ca_w_2_400_s_0_300 = 5.86e-05  mcm5m4l1_cc_w_2_400_s_0_300 = 9.20e-11  mcm5m4l1_cf_w_2_400_s_0_300 = 9.20e-12
+ mcm5m4l1_ca_w_2_400_s_0_360 = 5.86e-05  mcm5m4l1_cc_w_2_400_s_0_360 = 8.51e-11  mcm5m4l1_cf_w_2_400_s_0_360 = 1.07e-11
+ mcm5m4l1_ca_w_2_400_s_0_450 = 5.86e-05  mcm5m4l1_cc_w_2_400_s_0_450 = 7.59e-11  mcm5m4l1_cf_w_2_400_s_0_450 = 1.29e-11
+ mcm5m4l1_ca_w_2_400_s_0_600 = 5.86e-05  mcm5m4l1_cc_w_2_400_s_0_600 = 6.34e-11  mcm5m4l1_cf_w_2_400_s_0_600 = 1.64e-11
+ mcm5m4l1_ca_w_2_400_s_0_800 = 5.86e-05  mcm5m4l1_cc_w_2_400_s_0_800 = 5.06e-11  mcm5m4l1_cf_w_2_400_s_0_800 = 2.06e-11
+ mcm5m4l1_ca_w_2_400_s_1_000 = 5.86e-05  mcm5m4l1_cc_w_2_400_s_1_000 = 4.10e-11  mcm5m4l1_cf_w_2_400_s_1_000 = 2.44e-11
+ mcm5m4l1_ca_w_2_400_s_1_200 = 5.86e-05  mcm5m4l1_cc_w_2_400_s_1_200 = 3.37e-11  mcm5m4l1_cf_w_2_400_s_1_200 = 2.78e-11
+ mcm5m4l1_ca_w_2_400_s_2_100 = 5.86e-05  mcm5m4l1_cc_w_2_400_s_2_100 = 1.60e-11  mcm5m4l1_cf_w_2_400_s_2_100 = 3.87e-11
+ mcm5m4l1_ca_w_2_400_s_3_300 = 5.86e-05  mcm5m4l1_cc_w_2_400_s_3_300 = 6.82e-12  mcm5m4l1_cf_w_2_400_s_3_300 = 4.63e-11
+ mcm5m4l1_ca_w_2_400_s_9_000 = 5.86e-05  mcm5m4l1_cc_w_2_400_s_9_000 = 2.05e-13  mcm5m4l1_cf_w_2_400_s_9_000 = 5.25e-11
+ mcm5m4m1_ca_w_0_300_s_0_300 = 6.14e-05  mcm5m4m1_cc_w_0_300_s_0_300 = 8.11e-11  mcm5m4m1_cf_w_0_300_s_0_300 = 9.60e-12
+ mcm5m4m1_ca_w_0_300_s_0_360 = 6.14e-05  mcm5m4m1_cc_w_0_300_s_0_360 = 7.45e-11  mcm5m4m1_cf_w_0_300_s_0_360 = 1.12e-11
+ mcm5m4m1_ca_w_0_300_s_0_450 = 6.14e-05  mcm5m4m1_cc_w_0_300_s_0_450 = 6.62e-11  mcm5m4m1_cf_w_0_300_s_0_450 = 1.35e-11
+ mcm5m4m1_ca_w_0_300_s_0_600 = 6.14e-05  mcm5m4m1_cc_w_0_300_s_0_600 = 5.48e-11  mcm5m4m1_cf_w_0_300_s_0_600 = 1.72e-11
+ mcm5m4m1_ca_w_0_300_s_0_800 = 6.14e-05  mcm5m4m1_cc_w_0_300_s_0_800 = 4.32e-11  mcm5m4m1_cf_w_0_300_s_0_800 = 2.15e-11
+ mcm5m4m1_ca_w_0_300_s_1_000 = 6.14e-05  mcm5m4m1_cc_w_0_300_s_1_000 = 3.45e-11  mcm5m4m1_cf_w_0_300_s_1_000 = 2.54e-11
+ mcm5m4m1_ca_w_0_300_s_1_200 = 6.14e-05  mcm5m4m1_cc_w_0_300_s_1_200 = 2.79e-11  mcm5m4m1_cf_w_0_300_s_1_200 = 2.88e-11
+ mcm5m4m1_ca_w_0_300_s_2_100 = 6.14e-05  mcm5m4m1_cc_w_0_300_s_2_100 = 1.19e-11  mcm5m4m1_cf_w_0_300_s_2_100 = 3.94e-11
+ mcm5m4m1_ca_w_0_300_s_3_300 = 6.14e-05  mcm5m4m1_cc_w_0_300_s_3_300 = 4.41e-12  mcm5m4m1_cf_w_0_300_s_3_300 = 4.59e-11
+ mcm5m4m1_ca_w_0_300_s_9_000 = 6.14e-05  mcm5m4m1_cc_w_0_300_s_9_000 = 1.05e-13  mcm5m4m1_cf_w_0_300_s_9_000 = 5.01e-11
+ mcm5m4m1_ca_w_2_400_s_0_300 = 6.14e-05  mcm5m4m1_cc_w_2_400_s_0_300 = 8.98e-11  mcm5m4m1_cf_w_2_400_s_0_300 = 9.68e-12
+ mcm5m4m1_ca_w_2_400_s_0_360 = 6.14e-05  mcm5m4m1_cc_w_2_400_s_0_360 = 8.28e-11  mcm5m4m1_cf_w_2_400_s_0_360 = 1.13e-11
+ mcm5m4m1_ca_w_2_400_s_0_450 = 6.14e-05  mcm5m4m1_cc_w_2_400_s_0_450 = 7.37e-11  mcm5m4m1_cf_w_2_400_s_0_450 = 1.36e-11
+ mcm5m4m1_ca_w_2_400_s_0_600 = 6.14e-05  mcm5m4m1_cc_w_2_400_s_0_600 = 6.11e-11  mcm5m4m1_cf_w_2_400_s_0_600 = 1.72e-11
+ mcm5m4m1_ca_w_2_400_s_0_800 = 6.14e-05  mcm5m4m1_cc_w_2_400_s_0_800 = 4.83e-11  mcm5m4m1_cf_w_2_400_s_0_800 = 2.16e-11
+ mcm5m4m1_ca_w_2_400_s_1_000 = 6.14e-05  mcm5m4m1_cc_w_2_400_s_1_000 = 3.86e-11  mcm5m4m1_cf_w_2_400_s_1_000 = 2.56e-11
+ mcm5m4m1_ca_w_2_400_s_1_200 = 6.14e-05  mcm5m4m1_cc_w_2_400_s_1_200 = 3.14e-11  mcm5m4m1_cf_w_2_400_s_1_200 = 2.91e-11
+ mcm5m4m1_ca_w_2_400_s_2_100 = 6.14e-05  mcm5m4m1_cc_w_2_400_s_2_100 = 1.40e-11  mcm5m4m1_cf_w_2_400_s_2_100 = 4.04e-11
+ mcm5m4m1_ca_w_2_400_s_3_300 = 6.14e-05  mcm5m4m1_cc_w_2_400_s_3_300 = 5.31e-12  mcm5m4m1_cf_w_2_400_s_3_300 = 4.77e-11
+ mcm5m4m1_ca_w_2_400_s_9_000 = 6.14e-05  mcm5m4m1_cc_w_2_400_s_9_000 = 1.25e-13  mcm5m4m1_cf_w_2_400_s_9_000 = 5.27e-11
+ mcm5m4m2_ca_w_0_300_s_0_300 = 6.64e-05  mcm5m4m2_cc_w_0_300_s_0_300 = 7.98e-11  mcm5m4m2_cf_w_0_300_s_0_300 = 1.04e-11
+ mcm5m4m2_ca_w_0_300_s_0_360 = 6.64e-05  mcm5m4m2_cc_w_0_300_s_0_360 = 7.32e-11  mcm5m4m2_cf_w_0_300_s_0_360 = 1.21e-11
+ mcm5m4m2_ca_w_0_300_s_0_450 = 6.64e-05  mcm5m4m2_cc_w_0_300_s_0_450 = 6.47e-11  mcm5m4m2_cf_w_0_300_s_0_450 = 1.46e-11
+ mcm5m4m2_ca_w_0_300_s_0_600 = 6.64e-05  mcm5m4m2_cc_w_0_300_s_0_600 = 5.32e-11  mcm5m4m2_cf_w_0_300_s_0_600 = 1.86e-11
+ mcm5m4m2_ca_w_0_300_s_0_800 = 6.64e-05  mcm5m4m2_cc_w_0_300_s_0_800 = 4.13e-11  mcm5m4m2_cf_w_0_300_s_0_800 = 2.33e-11
+ mcm5m4m2_ca_w_0_300_s_1_000 = 6.64e-05  mcm5m4m2_cc_w_0_300_s_1_000 = 3.25e-11  mcm5m4m2_cf_w_0_300_s_1_000 = 2.75e-11
+ mcm5m4m2_ca_w_0_300_s_1_200 = 6.64e-05  mcm5m4m2_cc_w_0_300_s_1_200 = 2.58e-11  mcm5m4m2_cf_w_0_300_s_1_200 = 3.11e-11
+ mcm5m4m2_ca_w_0_300_s_2_100 = 6.64e-05  mcm5m4m2_cc_w_0_300_s_2_100 = 1.01e-11  mcm5m4m2_cf_w_0_300_s_2_100 = 4.20e-11
+ mcm5m4m2_ca_w_0_300_s_3_300 = 6.64e-05  mcm5m4m2_cc_w_0_300_s_3_300 = 3.24e-12  mcm5m4m2_cf_w_0_300_s_3_300 = 4.82e-11
+ mcm5m4m2_ca_w_0_300_s_9_000 = 6.64e-05  mcm5m4m2_cc_w_0_300_s_9_000 = 4.50e-14  mcm5m4m2_cf_w_0_300_s_9_000 = 5.13e-11
+ mcm5m4m2_ca_w_2_400_s_0_300 = 6.64e-05  mcm5m4m2_cc_w_2_400_s_0_300 = 8.65e-11  mcm5m4m2_cf_w_2_400_s_0_300 = 1.05e-11
+ mcm5m4m2_ca_w_2_400_s_0_360 = 6.64e-05  mcm5m4m2_cc_w_2_400_s_0_360 = 7.95e-11  mcm5m4m2_cf_w_2_400_s_0_360 = 1.22e-11
+ mcm5m4m2_ca_w_2_400_s_0_450 = 6.64e-05  mcm5m4m2_cc_w_2_400_s_0_450 = 7.03e-11  mcm5m4m2_cf_w_2_400_s_0_450 = 1.47e-11
+ mcm5m4m2_ca_w_2_400_s_0_600 = 6.64e-05  mcm5m4m2_cc_w_2_400_s_0_600 = 5.77e-11  mcm5m4m2_cf_w_2_400_s_0_600 = 1.87e-11
+ mcm5m4m2_ca_w_2_400_s_0_800 = 6.64e-05  mcm5m4m2_cc_w_2_400_s_0_800 = 4.49e-11  mcm5m4m2_cf_w_2_400_s_0_800 = 2.35e-11
+ mcm5m4m2_ca_w_2_400_s_1_000 = 6.64e-05  mcm5m4m2_cc_w_2_400_s_1_000 = 3.53e-11  mcm5m4m2_cf_w_2_400_s_1_000 = 2.78e-11
+ mcm5m4m2_ca_w_2_400_s_1_200 = 6.64e-05  mcm5m4m2_cc_w_2_400_s_1_200 = 2.82e-11  mcm5m4m2_cf_w_2_400_s_1_200 = 3.15e-11
+ mcm5m4m2_ca_w_2_400_s_2_100 = 6.64e-05  mcm5m4m2_cc_w_2_400_s_2_100 = 1.12e-11  mcm5m4m2_cf_w_2_400_s_2_100 = 4.31e-11
+ mcm5m4m2_ca_w_2_400_s_3_300 = 6.64e-05  mcm5m4m2_cc_w_2_400_s_3_300 = 3.63e-12  mcm5m4m2_cf_w_2_400_s_3_300 = 4.97e-11
+ mcm5m4m2_ca_w_2_400_s_9_000 = 6.64e-05  mcm5m4m2_cc_w_2_400_s_9_000 = 4.50e-14  mcm5m4m2_cf_w_2_400_s_9_000 = 5.33e-11
+ mcm5m4m3_ca_w_0_300_s_0_300 = 1.06e-04  mcm5m4m3_cc_w_0_300_s_0_300 = 7.20e-11  mcm5m4m3_cf_w_0_300_s_0_300 = 1.66e-11
+ mcm5m4m3_ca_w_0_300_s_0_360 = 1.06e-04  mcm5m4m3_cc_w_0_300_s_0_360 = 6.53e-11  mcm5m4m3_cf_w_0_300_s_0_360 = 1.92e-11
+ mcm5m4m3_ca_w_0_300_s_0_450 = 1.06e-04  mcm5m4m3_cc_w_0_300_s_0_450 = 5.64e-11  mcm5m4m3_cf_w_0_300_s_0_450 = 2.30e-11
+ mcm5m4m3_ca_w_0_300_s_0_600 = 1.06e-04  mcm5m4m3_cc_w_0_300_s_0_600 = 4.41e-11  mcm5m4m3_cf_w_0_300_s_0_600 = 2.87e-11
+ mcm5m4m3_ca_w_0_300_s_0_800 = 1.06e-04  mcm5m4m3_cc_w_0_300_s_0_800 = 3.21e-11  mcm5m4m3_cf_w_0_300_s_0_800 = 3.55e-11
+ mcm5m4m3_ca_w_0_300_s_1_000 = 1.06e-04  mcm5m4m3_cc_w_0_300_s_1_000 = 2.33e-11  mcm5m4m3_cf_w_0_300_s_1_000 = 4.11e-11
+ mcm5m4m3_ca_w_0_300_s_1_200 = 1.06e-04  mcm5m4m3_cc_w_0_300_s_1_200 = 1.70e-11  mcm5m4m3_cf_w_0_300_s_1_200 = 4.55e-11
+ mcm5m4m3_ca_w_0_300_s_2_100 = 1.06e-04  mcm5m4m3_cc_w_0_300_s_2_100 = 4.28e-12  mcm5m4m3_cf_w_0_300_s_2_100 = 5.62e-11
+ mcm5m4m3_ca_w_0_300_s_3_300 = 1.06e-04  mcm5m4m3_cc_w_0_300_s_3_300 = 7.20e-13  mcm5m4m3_cf_w_0_300_s_3_300 = 5.97e-11
+ mcm5m4m3_ca_w_0_300_s_9_000 = 1.06e-04  mcm5m4m3_cc_w_0_300_s_9_000 = 4.50e-14  mcm5m4m3_cf_w_0_300_s_9_000 = 6.05e-11
+ mcm5m4m3_ca_w_2_400_s_0_300 = 1.06e-04  mcm5m4m3_cc_w_2_400_s_0_300 = 7.38e-11  mcm5m4m3_cf_w_2_400_s_0_300 = 1.67e-11
+ mcm5m4m3_ca_w_2_400_s_0_360 = 1.06e-04  mcm5m4m3_cc_w_2_400_s_0_360 = 6.69e-11  mcm5m4m3_cf_w_2_400_s_0_360 = 1.93e-11
+ mcm5m4m3_ca_w_2_400_s_0_450 = 1.06e-04  mcm5m4m3_cc_w_2_400_s_0_450 = 5.76e-11  mcm5m4m3_cf_w_2_400_s_0_450 = 2.31e-11
+ mcm5m4m3_ca_w_2_400_s_0_600 = 1.06e-04  mcm5m4m3_cc_w_2_400_s_0_600 = 4.53e-11  mcm5m4m3_cf_w_2_400_s_0_600 = 2.89e-11
+ mcm5m4m3_ca_w_2_400_s_0_800 = 1.06e-04  mcm5m4m3_cc_w_2_400_s_0_800 = 3.29e-11  mcm5m4m3_cf_w_2_400_s_0_800 = 3.57e-11
+ mcm5m4m3_ca_w_2_400_s_1_000 = 1.06e-04  mcm5m4m3_cc_w_2_400_s_1_000 = 2.39e-11  mcm5m4m3_cf_w_2_400_s_1_000 = 4.14e-11
+ mcm5m4m3_ca_w_2_400_s_1_200 = 1.06e-04  mcm5m4m3_cc_w_2_400_s_1_200 = 1.74e-11  mcm5m4m3_cf_w_2_400_s_1_200 = 4.59e-11
+ mcm5m4m3_ca_w_2_400_s_2_100 = 1.06e-04  mcm5m4m3_cc_w_2_400_s_2_100 = 4.45e-12  mcm5m4m3_cf_w_2_400_s_2_100 = 5.68e-11
+ mcm5m4m3_ca_w_2_400_s_3_300 = 1.06e-04  mcm5m4m3_cc_w_2_400_s_3_300 = 7.50e-13  mcm5m4m3_cf_w_2_400_s_3_300 = 6.04e-11
+ mcm5m4m3_ca_w_2_400_s_9_000 = 1.06e-04  mcm5m4m3_cc_w_2_400_s_9_000 = 5.00e-14  mcm5m4m3_cf_w_2_400_s_9_000 = 6.12e-11
+ mcrdlm4f_ca_w_0_300_s_0_300 = 1.06e-05  mcrdlm4f_cc_w_0_300_s_0_300 = 9.24e-11  mcrdlm4f_cf_w_0_300_s_0_300 = 1.81e-12
+ mcrdlm4f_ca_w_0_300_s_0_360 = 1.06e-05  mcrdlm4f_cc_w_0_300_s_0_360 = 8.68e-11  mcrdlm4f_cf_w_0_300_s_0_360 = 2.13e-12
+ mcrdlm4f_ca_w_0_300_s_0_450 = 1.06e-05  mcrdlm4f_cc_w_0_300_s_0_450 = 7.89e-11  mcrdlm4f_cf_w_0_300_s_0_450 = 2.62e-12
+ mcrdlm4f_ca_w_0_300_s_0_600 = 1.06e-05  mcrdlm4f_cc_w_0_300_s_0_600 = 6.92e-11  mcrdlm4f_cf_w_0_300_s_0_600 = 3.42e-12
+ mcrdlm4f_ca_w_0_300_s_0_800 = 1.06e-05  mcrdlm4f_cc_w_0_300_s_0_800 = 5.94e-11  mcrdlm4f_cf_w_0_300_s_0_800 = 4.34e-12
+ mcrdlm4f_ca_w_0_300_s_1_000 = 1.06e-05  mcrdlm4f_cc_w_0_300_s_1_000 = 5.20e-11  mcrdlm4f_cf_w_0_300_s_1_000 = 5.32e-12
+ mcrdlm4f_ca_w_0_300_s_1_200 = 1.06e-05  mcrdlm4f_cc_w_0_300_s_1_200 = 4.62e-11  mcrdlm4f_cf_w_0_300_s_1_200 = 6.28e-12
+ mcrdlm4f_ca_w_0_300_s_2_100 = 1.06e-05  mcrdlm4f_cc_w_0_300_s_2_100 = 3.10e-11  mcrdlm4f_cf_w_0_300_s_2_100 = 1.05e-11
+ mcrdlm4f_ca_w_0_300_s_3_300 = 1.06e-05  mcrdlm4f_cc_w_0_300_s_3_300 = 2.12e-11  mcrdlm4f_cf_w_0_300_s_3_300 = 1.47e-11
+ mcrdlm4f_ca_w_0_300_s_9_000 = 1.06e-05  mcrdlm4f_cc_w_0_300_s_9_000 = 4.90e-12  mcrdlm4f_cf_w_0_300_s_9_000 = 2.60e-11
+ mcrdlm4f_ca_w_2_400_s_0_300 = 1.06e-05  mcrdlm4f_cc_w_2_400_s_0_300 = 1.18e-10  mcrdlm4f_cf_w_2_400_s_0_300 = 1.84e-12
+ mcrdlm4f_ca_w_2_400_s_0_360 = 1.06e-05  mcrdlm4f_cc_w_2_400_s_0_360 = 1.11e-10  mcrdlm4f_cf_w_2_400_s_0_360 = 2.15e-12
+ mcrdlm4f_ca_w_2_400_s_0_450 = 1.06e-05  mcrdlm4f_cc_w_2_400_s_0_450 = 1.02e-10  mcrdlm4f_cf_w_2_400_s_0_450 = 2.61e-12
+ mcrdlm4f_ca_w_2_400_s_0_600 = 1.06e-05  mcrdlm4f_cc_w_2_400_s_0_600 = 8.97e-11  mcrdlm4f_cf_w_2_400_s_0_600 = 3.38e-12
+ mcrdlm4f_ca_w_2_400_s_0_800 = 1.06e-05  mcrdlm4f_cc_w_2_400_s_0_800 = 7.71e-11  mcrdlm4f_cf_w_2_400_s_0_800 = 4.39e-12
+ mcrdlm4f_ca_w_2_400_s_1_000 = 1.06e-05  mcrdlm4f_cc_w_2_400_s_1_000 = 6.74e-11  mcrdlm4f_cf_w_2_400_s_1_000 = 5.38e-12
+ mcrdlm4f_ca_w_2_400_s_1_200 = 1.06e-05  mcrdlm4f_cc_w_2_400_s_1_200 = 6.00e-11  mcrdlm4f_cf_w_2_400_s_1_200 = 6.35e-12
+ mcrdlm4f_ca_w_2_400_s_2_100 = 1.06e-05  mcrdlm4f_cc_w_2_400_s_2_100 = 4.06e-11  mcrdlm4f_cf_w_2_400_s_2_100 = 1.05e-11
+ mcrdlm4f_ca_w_2_400_s_3_300 = 1.06e-05  mcrdlm4f_cc_w_2_400_s_3_300 = 2.76e-11  mcrdlm4f_cf_w_2_400_s_3_300 = 1.53e-11
+ mcrdlm4f_ca_w_2_400_s_9_000 = 1.06e-05  mcrdlm4f_cc_w_2_400_s_9_000 = 6.65e-12  mcrdlm4f_cf_w_2_400_s_9_000 = 2.87e-11
+ mcrdlm4d_ca_w_0_300_s_0_300 = 1.12e-05  mcrdlm4d_cc_w_0_300_s_0_300 = 9.22e-11  mcrdlm4d_cf_w_0_300_s_0_300 = 1.93e-12
+ mcrdlm4d_ca_w_0_300_s_0_360 = 1.12e-05  mcrdlm4d_cc_w_0_300_s_0_360 = 8.66e-11  mcrdlm4d_cf_w_0_300_s_0_360 = 2.27e-12
+ mcrdlm4d_ca_w_0_300_s_0_450 = 1.12e-05  mcrdlm4d_cc_w_0_300_s_0_450 = 7.87e-11  mcrdlm4d_cf_w_0_300_s_0_450 = 2.79e-12
+ mcrdlm4d_ca_w_0_300_s_0_600 = 1.12e-05  mcrdlm4d_cc_w_0_300_s_0_600 = 6.90e-11  mcrdlm4d_cf_w_0_300_s_0_600 = 3.64e-12
+ mcrdlm4d_ca_w_0_300_s_0_800 = 1.12e-05  mcrdlm4d_cc_w_0_300_s_0_800 = 5.92e-11  mcrdlm4d_cf_w_0_300_s_0_800 = 4.62e-12
+ mcrdlm4d_ca_w_0_300_s_1_000 = 1.12e-05  mcrdlm4d_cc_w_0_300_s_1_000 = 5.16e-11  mcrdlm4d_cf_w_0_300_s_1_000 = 5.65e-12
+ mcrdlm4d_ca_w_0_300_s_1_200 = 1.12e-05  mcrdlm4d_cc_w_0_300_s_1_200 = 4.58e-11  mcrdlm4d_cf_w_0_300_s_1_200 = 6.68e-12
+ mcrdlm4d_ca_w_0_300_s_2_100 = 1.12e-05  mcrdlm4d_cc_w_0_300_s_2_100 = 3.05e-11  mcrdlm4d_cf_w_0_300_s_2_100 = 1.11e-11
+ mcrdlm4d_ca_w_0_300_s_3_300 = 1.12e-05  mcrdlm4d_cc_w_0_300_s_3_300 = 2.06e-11  mcrdlm4d_cf_w_0_300_s_3_300 = 1.55e-11
+ mcrdlm4d_ca_w_0_300_s_9_000 = 1.12e-05  mcrdlm4d_cc_w_0_300_s_9_000 = 4.51e-12  mcrdlm4d_cf_w_0_300_s_9_000 = 2.69e-11
+ mcrdlm4d_ca_w_2_400_s_0_300 = 1.12e-05  mcrdlm4d_cc_w_2_400_s_0_300 = 1.17e-10  mcrdlm4d_cf_w_2_400_s_0_300 = 1.96e-12
+ mcrdlm4d_ca_w_2_400_s_0_360 = 1.12e-05  mcrdlm4d_cc_w_2_400_s_0_360 = 1.10e-10  mcrdlm4d_cf_w_2_400_s_0_360 = 2.29e-12
+ mcrdlm4d_ca_w_2_400_s_0_450 = 1.12e-05  mcrdlm4d_cc_w_2_400_s_0_450 = 1.01e-10  mcrdlm4d_cf_w_2_400_s_0_450 = 2.78e-12
+ mcrdlm4d_ca_w_2_400_s_0_600 = 1.12e-05  mcrdlm4d_cc_w_2_400_s_0_600 = 8.90e-11  mcrdlm4d_cf_w_2_400_s_0_600 = 3.60e-12
+ mcrdlm4d_ca_w_2_400_s_0_800 = 1.12e-05  mcrdlm4d_cc_w_2_400_s_0_800 = 7.65e-11  mcrdlm4d_cf_w_2_400_s_0_800 = 4.67e-12
+ mcrdlm4d_ca_w_2_400_s_1_000 = 1.12e-05  mcrdlm4d_cc_w_2_400_s_1_000 = 6.66e-11  mcrdlm4d_cf_w_2_400_s_1_000 = 5.72e-12
+ mcrdlm4d_ca_w_2_400_s_1_200 = 1.12e-05  mcrdlm4d_cc_w_2_400_s_1_200 = 5.93e-11  mcrdlm4d_cf_w_2_400_s_1_200 = 6.75e-12
+ mcrdlm4d_ca_w_2_400_s_2_100 = 1.12e-05  mcrdlm4d_cc_w_2_400_s_2_100 = 3.98e-11  mcrdlm4d_cf_w_2_400_s_2_100 = 1.11e-11
+ mcrdlm4d_ca_w_2_400_s_3_300 = 1.12e-05  mcrdlm4d_cc_w_2_400_s_3_300 = 2.67e-11  mcrdlm4d_cf_w_2_400_s_3_300 = 1.61e-11
+ mcrdlm4d_ca_w_2_400_s_9_000 = 1.12e-05  mcrdlm4d_cc_w_2_400_s_9_000 = 6.15e-12  mcrdlm4d_cf_w_2_400_s_9_000 = 2.97e-11
+ mcrdlm4p1_ca_w_0_300_s_0_300 = 1.17e-05  mcrdlm4p1_cc_w_0_300_s_0_300 = 9.21e-11  mcrdlm4p1_cf_w_0_300_s_0_300 = 2.01e-12
+ mcrdlm4p1_ca_w_0_300_s_0_360 = 1.17e-05  mcrdlm4p1_cc_w_0_300_s_0_360 = 8.65e-11  mcrdlm4p1_cf_w_0_300_s_0_360 = 2.36e-12
+ mcrdlm4p1_ca_w_0_300_s_0_450 = 1.17e-05  mcrdlm4p1_cc_w_0_300_s_0_450 = 7.86e-11  mcrdlm4p1_cf_w_0_300_s_0_450 = 2.90e-12
+ mcrdlm4p1_ca_w_0_300_s_0_600 = 1.17e-05  mcrdlm4p1_cc_w_0_300_s_0_600 = 6.88e-11  mcrdlm4p1_cf_w_0_300_s_0_600 = 3.78e-12
+ mcrdlm4p1_ca_w_0_300_s_0_800 = 1.17e-05  mcrdlm4p1_cc_w_0_300_s_0_800 = 5.89e-11  mcrdlm4p1_cf_w_0_300_s_0_800 = 4.79e-12
+ mcrdlm4p1_ca_w_0_300_s_1_000 = 1.17e-05  mcrdlm4p1_cc_w_0_300_s_1_000 = 5.13e-11  mcrdlm4p1_cf_w_0_300_s_1_000 = 5.87e-12
+ mcrdlm4p1_ca_w_0_300_s_1_200 = 1.17e-05  mcrdlm4p1_cc_w_0_300_s_1_200 = 4.55e-11  mcrdlm4p1_cf_w_0_300_s_1_200 = 6.93e-12
+ mcrdlm4p1_ca_w_0_300_s_2_100 = 1.17e-05  mcrdlm4p1_cc_w_0_300_s_2_100 = 3.02e-11  mcrdlm4p1_cf_w_0_300_s_2_100 = 1.15e-11
+ mcrdlm4p1_ca_w_0_300_s_3_300 = 1.17e-05  mcrdlm4p1_cc_w_0_300_s_3_300 = 2.02e-11  mcrdlm4p1_cf_w_0_300_s_3_300 = 1.60e-11
+ mcrdlm4p1_ca_w_0_300_s_9_000 = 1.17e-05  mcrdlm4p1_cc_w_0_300_s_9_000 = 4.30e-12  mcrdlm4p1_cf_w_0_300_s_9_000 = 2.74e-11
+ mcrdlm4p1_ca_w_2_400_s_0_300 = 1.17e-05  mcrdlm4p1_cc_w_2_400_s_0_300 = 1.17e-10  mcrdlm4p1_cf_w_2_400_s_0_300 = 2.04e-12
+ mcrdlm4p1_ca_w_2_400_s_0_360 = 1.17e-05  mcrdlm4p1_cc_w_2_400_s_0_360 = 1.10e-10  mcrdlm4p1_cf_w_2_400_s_0_360 = 2.38e-12
+ mcrdlm4p1_ca_w_2_400_s_0_450 = 1.17e-05  mcrdlm4p1_cc_w_2_400_s_0_450 = 1.01e-10  mcrdlm4p1_cf_w_2_400_s_0_450 = 2.90e-12
+ mcrdlm4p1_ca_w_2_400_s_0_600 = 1.17e-05  mcrdlm4p1_cc_w_2_400_s_0_600 = 8.86e-11  mcrdlm4p1_cf_w_2_400_s_0_600 = 3.74e-12
+ mcrdlm4p1_ca_w_2_400_s_0_800 = 1.17e-05  mcrdlm4p1_cc_w_2_400_s_0_800 = 7.60e-11  mcrdlm4p1_cf_w_2_400_s_0_800 = 4.85e-12
+ mcrdlm4p1_ca_w_2_400_s_1_000 = 1.17e-05  mcrdlm4p1_cc_w_2_400_s_1_000 = 6.62e-11  mcrdlm4p1_cf_w_2_400_s_1_000 = 5.94e-12
+ mcrdlm4p1_ca_w_2_400_s_1_200 = 1.17e-05  mcrdlm4p1_cc_w_2_400_s_1_200 = 5.88e-11  mcrdlm4p1_cf_w_2_400_s_1_200 = 7.00e-12
+ mcrdlm4p1_ca_w_2_400_s_2_100 = 1.17e-05  mcrdlm4p1_cc_w_2_400_s_2_100 = 3.93e-11  mcrdlm4p1_cf_w_2_400_s_2_100 = 1.15e-11
+ mcrdlm4p1_ca_w_2_400_s_3_300 = 1.17e-05  mcrdlm4p1_cc_w_2_400_s_3_300 = 2.62e-11  mcrdlm4p1_cf_w_2_400_s_3_300 = 1.67e-11
+ mcrdlm4p1_ca_w_2_400_s_9_000 = 1.17e-05  mcrdlm4p1_cc_w_2_400_s_9_000 = 5.86e-12  mcrdlm4p1_cf_w_2_400_s_9_000 = 3.03e-11
+ mcrdlm4l1_ca_w_0_300_s_0_300 = 1.32e-05  mcrdlm4l1_cc_w_0_300_s_0_300 = 9.17e-11  mcrdlm4l1_cf_w_0_300_s_0_300 = 2.26e-12
+ mcrdlm4l1_ca_w_0_300_s_0_360 = 1.32e-05  mcrdlm4l1_cc_w_0_300_s_0_360 = 8.60e-11  mcrdlm4l1_cf_w_0_300_s_0_360 = 2.65e-12
+ mcrdlm4l1_ca_w_0_300_s_0_450 = 1.32e-05  mcrdlm4l1_cc_w_0_300_s_0_450 = 7.82e-11  mcrdlm4l1_cf_w_0_300_s_0_450 = 3.26e-12
+ mcrdlm4l1_ca_w_0_300_s_0_600 = 1.32e-05  mcrdlm4l1_cc_w_0_300_s_0_600 = 6.83e-11  mcrdlm4l1_cf_w_0_300_s_0_600 = 4.24e-12
+ mcrdlm4l1_ca_w_0_300_s_0_800 = 1.32e-05  mcrdlm4l1_cc_w_0_300_s_0_800 = 5.85e-11  mcrdlm4l1_cf_w_0_300_s_0_800 = 5.39e-12
+ mcrdlm4l1_ca_w_0_300_s_1_000 = 1.32e-05  mcrdlm4l1_cc_w_0_300_s_1_000 = 5.06e-11  mcrdlm4l1_cf_w_0_300_s_1_000 = 6.57e-12
+ mcrdlm4l1_ca_w_0_300_s_1_200 = 1.32e-05  mcrdlm4l1_cc_w_0_300_s_1_200 = 4.48e-11  mcrdlm4l1_cf_w_0_300_s_1_200 = 7.73e-12
+ mcrdlm4l1_ca_w_0_300_s_2_100 = 1.32e-05  mcrdlm4l1_cc_w_0_300_s_2_100 = 2.91e-11  mcrdlm4l1_cf_w_0_300_s_2_100 = 1.27e-11
+ mcrdlm4l1_ca_w_0_300_s_3_300 = 1.32e-05  mcrdlm4l1_cc_w_0_300_s_3_300 = 1.91e-11  mcrdlm4l1_cf_w_0_300_s_3_300 = 1.76e-11
+ mcrdlm4l1_ca_w_0_300_s_9_000 = 1.32e-05  mcrdlm4l1_cc_w_0_300_s_9_000 = 3.69e-12  mcrdlm4l1_cf_w_0_300_s_9_000 = 2.90e-11
+ mcrdlm4l1_ca_w_2_400_s_0_300 = 1.32e-05  mcrdlm4l1_cc_w_2_400_s_0_300 = 1.15e-10  mcrdlm4l1_cf_w_2_400_s_0_300 = 2.28e-12
+ mcrdlm4l1_ca_w_2_400_s_0_360 = 1.32e-05  mcrdlm4l1_cc_w_2_400_s_0_360 = 1.09e-10  mcrdlm4l1_cf_w_2_400_s_0_360 = 2.66e-12
+ mcrdlm4l1_ca_w_2_400_s_0_450 = 1.32e-05  mcrdlm4l1_cc_w_2_400_s_0_450 = 9.95e-11  mcrdlm4l1_cf_w_2_400_s_0_450 = 3.24e-12
+ mcrdlm4l1_ca_w_2_400_s_0_600 = 1.32e-05  mcrdlm4l1_cc_w_2_400_s_0_600 = 8.72e-11  mcrdlm4l1_cf_w_2_400_s_0_600 = 4.18e-12
+ mcrdlm4l1_ca_w_2_400_s_0_800 = 1.32e-05  mcrdlm4l1_cc_w_2_400_s_0_800 = 7.46e-11  mcrdlm4l1_cf_w_2_400_s_0_800 = 5.43e-12
+ mcrdlm4l1_ca_w_2_400_s_1_000 = 1.32e-05  mcrdlm4l1_cc_w_2_400_s_1_000 = 6.48e-11  mcrdlm4l1_cf_w_2_400_s_1_000 = 6.63e-12
+ mcrdlm4l1_ca_w_2_400_s_1_200 = 1.32e-05  mcrdlm4l1_cc_w_2_400_s_1_200 = 5.74e-11  mcrdlm4l1_cf_w_2_400_s_1_200 = 7.81e-12
+ mcrdlm4l1_ca_w_2_400_s_2_100 = 1.32e-05  mcrdlm4l1_cc_w_2_400_s_2_100 = 3.78e-11  mcrdlm4l1_cf_w_2_400_s_2_100 = 1.28e-11
+ mcrdlm4l1_ca_w_2_400_s_3_300 = 1.32e-05  mcrdlm4l1_cc_w_2_400_s_3_300 = 2.48e-11  mcrdlm4l1_cf_w_2_400_s_3_300 = 1.83e-11
+ mcrdlm4l1_ca_w_2_400_s_9_000 = 1.32e-05  mcrdlm4l1_cc_w_2_400_s_9_000 = 5.06e-12  mcrdlm4l1_cf_w_2_400_s_9_000 = 3.21e-11
+ mcrdlm4m1_ca_w_0_300_s_0_300 = 1.60e-05  mcrdlm4m1_cc_w_0_300_s_0_300 = 9.09e-11  mcrdlm4m1_cf_w_0_300_s_0_300 = 2.73e-12
+ mcrdlm4m1_ca_w_0_300_s_0_360 = 1.60e-05  mcrdlm4m1_cc_w_0_300_s_0_360 = 8.53e-11  mcrdlm4m1_cf_w_0_300_s_0_360 = 3.20e-12
+ mcrdlm4m1_ca_w_0_300_s_0_450 = 1.60e-05  mcrdlm4m1_cc_w_0_300_s_0_450 = 7.75e-11  mcrdlm4m1_cf_w_0_300_s_0_450 = 3.93e-12
+ mcrdlm4m1_ca_w_0_300_s_0_600 = 1.60e-05  mcrdlm4m1_cc_w_0_300_s_0_600 = 6.73e-11  mcrdlm4m1_cf_w_0_300_s_0_600 = 5.10e-12
+ mcrdlm4m1_ca_w_0_300_s_0_800 = 1.60e-05  mcrdlm4m1_cc_w_0_300_s_0_800 = 5.73e-11  mcrdlm4m1_cf_w_0_300_s_0_800 = 6.49e-12
+ mcrdlm4m1_ca_w_0_300_s_1_000 = 1.60e-05  mcrdlm4m1_cc_w_0_300_s_1_000 = 4.94e-11  mcrdlm4m1_cf_w_0_300_s_1_000 = 7.87e-12
+ mcrdlm4m1_ca_w_0_300_s_1_200 = 1.60e-05  mcrdlm4m1_cc_w_0_300_s_1_200 = 4.33e-11  mcrdlm4m1_cf_w_0_300_s_1_200 = 9.24e-12
+ mcrdlm4m1_ca_w_0_300_s_2_100 = 1.60e-05  mcrdlm4m1_cc_w_0_300_s_2_100 = 2.74e-11  mcrdlm4m1_cf_w_0_300_s_2_100 = 1.50e-11
+ mcrdlm4m1_ca_w_0_300_s_3_300 = 1.60e-05  mcrdlm4m1_cc_w_0_300_s_3_300 = 1.73e-11  mcrdlm4m1_cf_w_0_300_s_3_300 = 2.04e-11
+ mcrdlm4m1_ca_w_0_300_s_9_000 = 1.60e-05  mcrdlm4m1_cc_w_0_300_s_9_000 = 2.88e-12  mcrdlm4m1_cf_w_0_300_s_9_000 = 3.17e-11
+ mcrdlm4m1_ca_w_2_400_s_0_300 = 1.60e-05  mcrdlm4m1_cc_w_2_400_s_0_300 = 1.14e-10  mcrdlm4m1_cf_w_2_400_s_0_300 = 2.75e-12
+ mcrdlm4m1_ca_w_2_400_s_0_360 = 1.60e-05  mcrdlm4m1_cc_w_2_400_s_0_360 = 1.06e-10  mcrdlm4m1_cf_w_2_400_s_0_360 = 3.21e-12
+ mcrdlm4m1_ca_w_2_400_s_0_450 = 1.60e-05  mcrdlm4m1_cc_w_2_400_s_0_450 = 9.72e-11  mcrdlm4m1_cf_w_2_400_s_0_450 = 3.90e-12
+ mcrdlm4m1_ca_w_2_400_s_0_600 = 1.60e-05  mcrdlm4m1_cc_w_2_400_s_0_600 = 8.49e-11  mcrdlm4m1_cf_w_2_400_s_0_600 = 5.04e-12
+ mcrdlm4m1_ca_w_2_400_s_0_800 = 1.60e-05  mcrdlm4m1_cc_w_2_400_s_0_800 = 7.22e-11  mcrdlm4m1_cf_w_2_400_s_0_800 = 6.52e-12
+ mcrdlm4m1_ca_w_2_400_s_1_000 = 1.60e-05  mcrdlm4m1_cc_w_2_400_s_1_000 = 6.25e-11  mcrdlm4m1_cf_w_2_400_s_1_000 = 7.97e-12
+ mcrdlm4m1_ca_w_2_400_s_1_200 = 1.60e-05  mcrdlm4m1_cc_w_2_400_s_1_200 = 5.50e-11  mcrdlm4m1_cf_w_2_400_s_1_200 = 9.35e-12
+ mcrdlm4m1_ca_w_2_400_s_2_100 = 1.60e-05  mcrdlm4m1_cc_w_2_400_s_2_100 = 3.53e-11  mcrdlm4m1_cf_w_2_400_s_2_100 = 1.51e-11
+ mcrdlm4m1_ca_w_2_400_s_3_300 = 1.60e-05  mcrdlm4m1_cc_w_2_400_s_3_300 = 2.25e-11  mcrdlm4m1_cf_w_2_400_s_3_300 = 2.13e-11
+ mcrdlm4m1_ca_w_2_400_s_9_000 = 1.60e-05  mcrdlm4m1_cc_w_2_400_s_9_000 = 4.02e-12  mcrdlm4m1_cf_w_2_400_s_9_000 = 3.51e-11
+ mcrdlm4m2_ca_w_0_300_s_0_300 = 2.10e-05  mcrdlm4m2_cc_w_0_300_s_0_300 = 8.94e-11  mcrdlm4m2_cf_w_0_300_s_0_300 = 3.56e-12
+ mcrdlm4m2_ca_w_0_300_s_0_360 = 2.10e-05  mcrdlm4m2_cc_w_0_300_s_0_360 = 8.40e-11  mcrdlm4m2_cf_w_0_300_s_0_360 = 4.16e-12
+ mcrdlm4m2_ca_w_0_300_s_0_450 = 2.10e-05  mcrdlm4m2_cc_w_0_300_s_0_450 = 7.61e-11  mcrdlm4m2_cf_w_0_300_s_0_450 = 5.08e-12
+ mcrdlm4m2_ca_w_0_300_s_0_600 = 2.10e-05  mcrdlm4m2_cc_w_0_300_s_0_600 = 6.57e-11  mcrdlm4m2_cf_w_0_300_s_0_600 = 6.57e-12
+ mcrdlm4m2_ca_w_0_300_s_0_800 = 2.10e-05  mcrdlm4m2_cc_w_0_300_s_0_800 = 5.54e-11  mcrdlm4m2_cf_w_0_300_s_0_800 = 8.35e-12
+ mcrdlm4m2_ca_w_0_300_s_1_000 = 2.10e-05  mcrdlm4m2_cc_w_0_300_s_1_000 = 4.73e-11  mcrdlm4m2_cf_w_0_300_s_1_000 = 1.01e-11
+ mcrdlm4m2_ca_w_0_300_s_1_200 = 2.10e-05  mcrdlm4m2_cc_w_0_300_s_1_200 = 4.11e-11  mcrdlm4m2_cf_w_0_300_s_1_200 = 1.18e-11
+ mcrdlm4m2_ca_w_0_300_s_2_100 = 2.10e-05  mcrdlm4m2_cc_w_0_300_s_2_100 = 2.49e-11  mcrdlm4m2_cf_w_0_300_s_2_100 = 1.86e-11
+ mcrdlm4m2_ca_w_0_300_s_3_300 = 2.10e-05  mcrdlm4m2_cc_w_0_300_s_3_300 = 1.49e-11  mcrdlm4m2_cf_w_0_300_s_3_300 = 2.47e-11
+ mcrdlm4m2_ca_w_0_300_s_9_000 = 2.10e-05  mcrdlm4m2_cc_w_0_300_s_9_000 = 2.04e-12  mcrdlm4m2_cf_w_0_300_s_9_000 = 3.54e-11
+ mcrdlm4m2_ca_w_2_400_s_0_300 = 2.10e-05  mcrdlm4m2_cc_w_2_400_s_0_300 = 1.10e-10  mcrdlm4m2_cf_w_2_400_s_0_300 = 3.58e-12
+ mcrdlm4m2_ca_w_2_400_s_0_360 = 2.10e-05  mcrdlm4m2_cc_w_2_400_s_0_360 = 1.03e-10  mcrdlm4m2_cf_w_2_400_s_0_360 = 4.18e-12
+ mcrdlm4m2_ca_w_2_400_s_0_450 = 2.10e-05  mcrdlm4m2_cc_w_2_400_s_0_450 = 9.38e-11  mcrdlm4m2_cf_w_2_400_s_0_450 = 5.07e-12
+ mcrdlm4m2_ca_w_2_400_s_0_600 = 2.10e-05  mcrdlm4m2_cc_w_2_400_s_0_600 = 8.15e-11  mcrdlm4m2_cf_w_2_400_s_0_600 = 6.52e-12
+ mcrdlm4m2_ca_w_2_400_s_0_800 = 2.10e-05  mcrdlm4m2_cc_w_2_400_s_0_800 = 6.88e-11  mcrdlm4m2_cf_w_2_400_s_0_800 = 8.40e-12
+ mcrdlm4m2_ca_w_2_400_s_1_000 = 2.10e-05  mcrdlm4m2_cc_w_2_400_s_1_000 = 5.91e-11  mcrdlm4m2_cf_w_2_400_s_1_000 = 1.02e-11
+ mcrdlm4m2_ca_w_2_400_s_1_200 = 2.10e-05  mcrdlm4m2_cc_w_2_400_s_1_200 = 5.17e-11  mcrdlm4m2_cf_w_2_400_s_1_200 = 1.19e-11
+ mcrdlm4m2_ca_w_2_400_s_2_100 = 2.10e-05  mcrdlm4m2_cc_w_2_400_s_2_100 = 3.21e-11  mcrdlm4m2_cf_w_2_400_s_2_100 = 1.88e-11
+ mcrdlm4m2_ca_w_2_400_s_3_300 = 2.10e-05  mcrdlm4m2_cc_w_2_400_s_3_300 = 1.96e-11  mcrdlm4m2_cf_w_2_400_s_3_300 = 2.58e-11
+ mcrdlm4m2_ca_w_2_400_s_9_000 = 2.10e-05  mcrdlm4m2_cc_w_2_400_s_9_000 = 2.96e-12  mcrdlm4m2_cf_w_2_400_s_9_000 = 3.91e-11
+ mcrdlm4m3_ca_w_0_300_s_0_300 = 6.09e-05  mcrdlm4m3_cc_w_0_300_s_0_300 = 8.16e-11  mcrdlm4m3_cf_w_0_300_s_0_300 = 9.73e-12
+ mcrdlm4m3_ca_w_0_300_s_0_360 = 6.09e-05  mcrdlm4m3_cc_w_0_300_s_0_360 = 7.59e-11  mcrdlm4m3_cf_w_0_300_s_0_360 = 1.12e-11
+ mcrdlm4m3_ca_w_0_300_s_0_450 = 6.09e-05  mcrdlm4m3_cc_w_0_300_s_0_450 = 6.75e-11  mcrdlm4m3_cf_w_0_300_s_0_450 = 1.35e-11
+ mcrdlm4m3_ca_w_0_300_s_0_600 = 6.09e-05  mcrdlm4m3_cc_w_0_300_s_0_600 = 5.66e-11  mcrdlm4m3_cf_w_0_300_s_0_600 = 1.69e-11
+ mcrdlm4m3_ca_w_0_300_s_0_800 = 6.09e-05  mcrdlm4m3_cc_w_0_300_s_0_800 = 4.58e-11  mcrdlm4m3_cf_w_0_300_s_0_800 = 2.08e-11
+ mcrdlm4m3_ca_w_0_300_s_1_000 = 6.09e-05  mcrdlm4m3_cc_w_0_300_s_1_000 = 3.76e-11  mcrdlm4m3_cf_w_0_300_s_1_000 = 2.44e-11
+ mcrdlm4m3_ca_w_0_300_s_1_200 = 6.09e-05  mcrdlm4m3_cc_w_0_300_s_1_200 = 3.14e-11  mcrdlm4m3_cf_w_0_300_s_1_200 = 2.75e-11
+ mcrdlm4m3_ca_w_0_300_s_2_100 = 6.09e-05  mcrdlm4m3_cc_w_0_300_s_2_100 = 1.58e-11  mcrdlm4m3_cf_w_0_300_s_2_100 = 3.78e-11
+ mcrdlm4m3_ca_w_0_300_s_3_300 = 6.09e-05  mcrdlm4m3_cc_w_0_300_s_3_300 = 8.00e-12  mcrdlm4m3_cf_w_0_300_s_3_300 = 4.43e-11
+ mcrdlm4m3_ca_w_0_300_s_9_000 = 6.09e-05  mcrdlm4m3_cc_w_0_300_s_9_000 = 7.20e-13  mcrdlm4m3_cf_w_0_300_s_9_000 = 5.11e-11
+ mcrdlm4m3_ca_w_2_400_s_0_300 = 6.09e-05  mcrdlm4m3_cc_w_2_400_s_0_300 = 9.75e-11  mcrdlm4m3_cf_w_2_400_s_0_300 = 9.75e-12
+ mcrdlm4m3_ca_w_2_400_s_0_360 = 6.09e-05  mcrdlm4m3_cc_w_2_400_s_0_360 = 9.06e-11  mcrdlm4m3_cf_w_2_400_s_0_360 = 1.13e-11
+ mcrdlm4m3_ca_w_2_400_s_0_450 = 6.09e-05  mcrdlm4m3_cc_w_2_400_s_0_450 = 8.14e-11  mcrdlm4m3_cf_w_2_400_s_0_450 = 1.35e-11
+ mcrdlm4m3_ca_w_2_400_s_0_600 = 6.09e-05  mcrdlm4m3_cc_w_2_400_s_0_600 = 6.91e-11  mcrdlm4m3_cf_w_2_400_s_0_600 = 1.69e-11
+ mcrdlm4m3_ca_w_2_400_s_0_800 = 6.09e-05  mcrdlm4m3_cc_w_2_400_s_0_800 = 5.66e-11  mcrdlm4m3_cf_w_2_400_s_0_800 = 2.09e-11
+ mcrdlm4m3_ca_w_2_400_s_1_000 = 6.09e-05  mcrdlm4m3_cc_w_2_400_s_1_000 = 4.72e-11  mcrdlm4m3_cf_w_2_400_s_1_000 = 2.46e-11
+ mcrdlm4m3_ca_w_2_400_s_1_200 = 6.09e-05  mcrdlm4m3_cc_w_2_400_s_1_200 = 4.01e-11  mcrdlm4m3_cf_w_2_400_s_1_200 = 2.78e-11
+ mcrdlm4m3_ca_w_2_400_s_2_100 = 6.09e-05  mcrdlm4m3_cc_w_2_400_s_2_100 = 2.23e-11  mcrdlm4m3_cf_w_2_400_s_2_100 = 3.83e-11
+ mcrdlm4m3_ca_w_2_400_s_3_300 = 6.09e-05  mcrdlm4m3_cc_w_2_400_s_3_300 = 1.20e-11  mcrdlm4m3_cf_w_2_400_s_3_300 = 4.63e-11
+ mcrdlm4m3_ca_w_2_400_s_9_000 = 6.09e-05  mcrdlm4m3_cc_w_2_400_s_9_000 = 1.24e-12  mcrdlm4m3_cf_w_2_400_s_9_000 = 5.62e-11
+ mcrdlm5f_ca_w_1_600_s_1_600 = 9.86e-06  mcrdlm5f_cc_w_1_600_s_1_600 = 5.94e-11  mcrdlm5f_cf_w_1_600_s_1_600 = 8.05e-12
+ mcrdlm5f_ca_w_1_600_s_1_700 = 9.86e-06  mcrdlm5f_cc_w_1_600_s_1_700 = 5.64e-11  mcrdlm5f_cf_w_1_600_s_1_700 = 8.49e-12
+ mcrdlm5f_ca_w_1_600_s_1_900 = 9.86e-06  mcrdlm5f_cc_w_1_600_s_1_900 = 5.14e-11  mcrdlm5f_cf_w_1_600_s_1_900 = 9.36e-12
+ mcrdlm5f_ca_w_1_600_s_2_000 = 9.86e-06  mcrdlm5f_cc_w_1_600_s_2_000 = 4.92e-11  mcrdlm5f_cf_w_1_600_s_2_000 = 9.78e-12
+ mcrdlm5f_ca_w_1_600_s_2_400 = 9.86e-06  mcrdlm5f_cc_w_1_600_s_2_400 = 4.21e-11  mcrdlm5f_cf_w_1_600_s_2_400 = 1.15e-11
+ mcrdlm5f_ca_w_1_600_s_2_800 = 9.86e-06  mcrdlm5f_cc_w_1_600_s_2_800 = 3.65e-11  mcrdlm5f_cf_w_1_600_s_2_800 = 1.31e-11
+ mcrdlm5f_ca_w_1_600_s_3_200 = 9.86e-06  mcrdlm5f_cc_w_1_600_s_3_200 = 3.21e-11  mcrdlm5f_cf_w_1_600_s_3_200 = 1.46e-11
+ mcrdlm5f_ca_w_1_600_s_4_800 = 9.86e-06  mcrdlm5f_cc_w_1_600_s_4_800 = 2.04e-11  mcrdlm5f_cf_w_1_600_s_4_800 = 2.00e-11
+ mcrdlm5f_ca_w_1_600_s_10_000 = 9.86e-06  mcrdlm5f_cc_w_1_600_s_10_000 = 5.89e-12  mcrdlm5f_cf_w_1_600_s_10_000 = 3.02e-11
+ mcrdlm5f_ca_w_1_600_s_12_000 = 9.86e-06  mcrdlm5f_cc_w_1_600_s_12_000 = 3.74e-12  mcrdlm5f_cf_w_1_600_s_12_000 = 3.20e-11
+ mcrdlm5f_ca_w_4_000_s_1_600 = 9.86e-06  mcrdlm5f_cc_w_4_000_s_1_600 = 6.35e-11  mcrdlm5f_cf_w_4_000_s_1_600 = 8.05e-12
+ mcrdlm5f_ca_w_4_000_s_1_700 = 9.86e-06  mcrdlm5f_cc_w_4_000_s_1_700 = 6.05e-11  mcrdlm5f_cf_w_4_000_s_1_700 = 8.50e-12
+ mcrdlm5f_ca_w_4_000_s_1_900 = 9.86e-06  mcrdlm5f_cc_w_4_000_s_1_900 = 5.52e-11  mcrdlm5f_cf_w_4_000_s_1_900 = 9.37e-12
+ mcrdlm5f_ca_w_4_000_s_2_000 = 9.86e-06  mcrdlm5f_cc_w_4_000_s_2_000 = 5.28e-11  mcrdlm5f_cf_w_4_000_s_2_000 = 9.82e-12
+ mcrdlm5f_ca_w_4_000_s_2_400 = 9.86e-06  mcrdlm5f_cc_w_4_000_s_2_400 = 4.50e-11  mcrdlm5f_cf_w_4_000_s_2_400 = 1.15e-11
+ mcrdlm5f_ca_w_4_000_s_2_800 = 9.86e-06  mcrdlm5f_cc_w_4_000_s_2_800 = 3.91e-11  mcrdlm5f_cf_w_4_000_s_2_800 = 1.31e-11
+ mcrdlm5f_ca_w_4_000_s_3_200 = 9.86e-06  mcrdlm5f_cc_w_4_000_s_3_200 = 3.44e-11  mcrdlm5f_cf_w_4_000_s_3_200 = 1.47e-11
+ mcrdlm5f_ca_w_4_000_s_4_800 = 9.86e-06  mcrdlm5f_cc_w_4_000_s_4_800 = 2.19e-11  mcrdlm5f_cf_w_4_000_s_4_800 = 2.02e-11
+ mcrdlm5f_ca_w_4_000_s_10_000 = 9.86e-06  mcrdlm5f_cc_w_4_000_s_10_000 = 6.41e-12  mcrdlm5f_cf_w_4_000_s_10_000 = 3.09e-11
+ mcrdlm5f_ca_w_4_000_s_12_000 = 9.86e-06  mcrdlm5f_cc_w_4_000_s_12_000 = 4.09e-12  mcrdlm5f_cf_w_4_000_s_12_000 = 3.29e-11
+ mcrdlm5d_ca_w_1_600_s_1_600 = 1.03e-05  mcrdlm5d_cc_w_1_600_s_1_600 = 5.90e-11  mcrdlm5d_cf_w_1_600_s_1_600 = 8.36e-12
+ mcrdlm5d_ca_w_1_600_s_1_700 = 1.03e-05  mcrdlm5d_cc_w_1_600_s_1_700 = 5.60e-11  mcrdlm5d_cf_w_1_600_s_1_700 = 8.83e-12
+ mcrdlm5d_ca_w_1_600_s_1_900 = 1.03e-05  mcrdlm5d_cc_w_1_600_s_1_900 = 5.10e-11  mcrdlm5d_cf_w_1_600_s_1_900 = 9.72e-12
+ mcrdlm5d_ca_w_1_600_s_2_000 = 1.03e-05  mcrdlm5d_cc_w_1_600_s_2_000 = 4.88e-11  mcrdlm5d_cf_w_1_600_s_2_000 = 1.02e-11
+ mcrdlm5d_ca_w_1_600_s_2_400 = 1.03e-05  mcrdlm5d_cc_w_1_600_s_2_400 = 4.15e-11  mcrdlm5d_cf_w_1_600_s_2_400 = 1.19e-11
+ mcrdlm5d_ca_w_1_600_s_2_800 = 1.03e-05  mcrdlm5d_cc_w_1_600_s_2_800 = 3.60e-11  mcrdlm5d_cf_w_1_600_s_2_800 = 1.36e-11
+ mcrdlm5d_ca_w_1_600_s_3_200 = 1.03e-05  mcrdlm5d_cc_w_1_600_s_3_200 = 3.16e-11  mcrdlm5d_cf_w_1_600_s_3_200 = 1.51e-11
+ mcrdlm5d_ca_w_1_600_s_4_800 = 1.03e-05  mcrdlm5d_cc_w_1_600_s_4_800 = 1.99e-11  mcrdlm5d_cf_w_1_600_s_4_800 = 2.06e-11
+ mcrdlm5d_ca_w_1_600_s_10_000 = 1.03e-05  mcrdlm5d_cc_w_1_600_s_10_000 = 5.53e-12  mcrdlm5d_cf_w_1_600_s_10_000 = 3.08e-11
+ mcrdlm5d_ca_w_1_600_s_12_000 = 1.03e-05  mcrdlm5d_cc_w_1_600_s_12_000 = 3.46e-12  mcrdlm5d_cf_w_1_600_s_12_000 = 3.27e-11
+ mcrdlm5d_ca_w_4_000_s_1_600 = 1.03e-05  mcrdlm5d_cc_w_4_000_s_1_600 = 6.29e-11  mcrdlm5d_cf_w_4_000_s_1_600 = 8.36e-12
+ mcrdlm5d_ca_w_4_000_s_1_700 = 1.03e-05  mcrdlm5d_cc_w_4_000_s_1_700 = 5.98e-11  mcrdlm5d_cf_w_4_000_s_1_700 = 8.83e-12
+ mcrdlm5d_ca_w_4_000_s_1_900 = 1.03e-05  mcrdlm5d_cc_w_4_000_s_1_900 = 5.45e-11  mcrdlm5d_cf_w_4_000_s_1_900 = 9.74e-12
+ mcrdlm5d_ca_w_4_000_s_2_000 = 1.03e-05  mcrdlm5d_cc_w_4_000_s_2_000 = 5.21e-11  mcrdlm5d_cf_w_4_000_s_2_000 = 1.02e-11
+ mcrdlm5d_ca_w_4_000_s_2_400 = 1.03e-05  mcrdlm5d_cc_w_4_000_s_2_400 = 4.44e-11  mcrdlm5d_cf_w_4_000_s_2_400 = 1.19e-11
+ mcrdlm5d_ca_w_4_000_s_2_800 = 1.03e-05  mcrdlm5d_cc_w_4_000_s_2_800 = 3.84e-11  mcrdlm5d_cf_w_4_000_s_2_800 = 1.36e-11
+ mcrdlm5d_ca_w_4_000_s_3_200 = 1.03e-05  mcrdlm5d_cc_w_4_000_s_3_200 = 3.37e-11  mcrdlm5d_cf_w_4_000_s_3_200 = 1.52e-11
+ mcrdlm5d_ca_w_4_000_s_4_800 = 1.03e-05  mcrdlm5d_cc_w_4_000_s_4_800 = 2.14e-11  mcrdlm5d_cf_w_4_000_s_4_800 = 2.08e-11
+ mcrdlm5d_ca_w_4_000_s_10_000 = 1.03e-05  mcrdlm5d_cc_w_4_000_s_10_000 = 5.99e-12  mcrdlm5d_cf_w_4_000_s_10_000 = 3.16e-11
+ mcrdlm5d_ca_w_4_000_s_12_000 = 1.03e-05  mcrdlm5d_cc_w_4_000_s_12_000 = 3.78e-12  mcrdlm5d_cf_w_4_000_s_12_000 = 3.36e-11
+ mcrdlm5p1_ca_w_1_600_s_1_600 = 1.05e-05  mcrdlm5p1_cc_w_1_600_s_1_600 = 5.87e-11  mcrdlm5p1_cf_w_1_600_s_1_600 = 8.56e-12
+ mcrdlm5p1_ca_w_1_600_s_1_700 = 1.05e-05  mcrdlm5p1_cc_w_1_600_s_1_700 = 5.57e-11  mcrdlm5p1_cf_w_1_600_s_1_700 = 9.02e-12
+ mcrdlm5p1_ca_w_1_600_s_1_900 = 1.05e-05  mcrdlm5p1_cc_w_1_600_s_1_900 = 5.07e-11  mcrdlm5p1_cf_w_1_600_s_1_900 = 9.95e-12
+ mcrdlm5p1_ca_w_1_600_s_2_000 = 1.05e-05  mcrdlm5p1_cc_w_1_600_s_2_000 = 4.85e-11  mcrdlm5p1_cf_w_1_600_s_2_000 = 1.04e-11
+ mcrdlm5p1_ca_w_1_600_s_2_400 = 1.05e-05  mcrdlm5p1_cc_w_1_600_s_2_400 = 4.12e-11  mcrdlm5p1_cf_w_1_600_s_2_400 = 1.22e-11
+ mcrdlm5p1_ca_w_1_600_s_2_800 = 1.05e-05  mcrdlm5p1_cc_w_1_600_s_2_800 = 3.57e-11  mcrdlm5p1_cf_w_1_600_s_2_800 = 1.39e-11
+ mcrdlm5p1_ca_w_1_600_s_3_200 = 1.05e-05  mcrdlm5p1_cc_w_1_600_s_3_200 = 3.13e-11  mcrdlm5p1_cf_w_1_600_s_3_200 = 1.55e-11
+ mcrdlm5p1_ca_w_1_600_s_4_800 = 1.05e-05  mcrdlm5p1_cc_w_1_600_s_4_800 = 1.96e-11  mcrdlm5p1_cf_w_1_600_s_4_800 = 2.11e-11
+ mcrdlm5p1_ca_w_1_600_s_10_000 = 1.05e-05  mcrdlm5p1_cc_w_1_600_s_10_000 = 5.31e-12  mcrdlm5p1_cf_w_1_600_s_10_000 = 3.13e-11
+ mcrdlm5p1_ca_w_1_600_s_12_000 = 1.05e-05  mcrdlm5p1_cc_w_1_600_s_12_000 = 3.29e-12  mcrdlm5p1_cf_w_1_600_s_12_000 = 3.31e-11
+ mcrdlm5p1_ca_w_4_000_s_1_600 = 1.05e-05  mcrdlm5p1_cc_w_4_000_s_1_600 = 6.25e-11  mcrdlm5p1_cf_w_4_000_s_1_600 = 8.56e-12
+ mcrdlm5p1_ca_w_4_000_s_1_700 = 1.05e-05  mcrdlm5p1_cc_w_4_000_s_1_700 = 5.94e-11  mcrdlm5p1_cf_w_4_000_s_1_700 = 9.04e-12
+ mcrdlm5p1_ca_w_4_000_s_1_900 = 1.05e-05  mcrdlm5p1_cc_w_4_000_s_1_900 = 5.40e-11  mcrdlm5p1_cf_w_4_000_s_1_900 = 9.97e-12
+ mcrdlm5p1_ca_w_4_000_s_2_000 = 1.05e-05  mcrdlm5p1_cc_w_4_000_s_2_000 = 5.17e-11  mcrdlm5p1_cf_w_4_000_s_2_000 = 1.04e-11
+ mcrdlm5p1_ca_w_4_000_s_2_400 = 1.05e-05  mcrdlm5p1_cc_w_4_000_s_2_400 = 4.40e-11  mcrdlm5p1_cf_w_4_000_s_2_400 = 1.22e-11
+ mcrdlm5p1_ca_w_4_000_s_2_800 = 1.05e-05  mcrdlm5p1_cc_w_4_000_s_2_800 = 3.81e-11  mcrdlm5p1_cf_w_4_000_s_2_800 = 1.39e-11
+ mcrdlm5p1_ca_w_4_000_s_3_200 = 1.05e-05  mcrdlm5p1_cc_w_4_000_s_3_200 = 3.34e-11  mcrdlm5p1_cf_w_4_000_s_3_200 = 1.56e-11
+ mcrdlm5p1_ca_w_4_000_s_4_800 = 1.05e-05  mcrdlm5p1_cc_w_4_000_s_4_800 = 2.10e-11  mcrdlm5p1_cf_w_4_000_s_4_800 = 2.13e-11
+ mcrdlm5p1_ca_w_4_000_s_10_000 = 1.05e-05  mcrdlm5p1_cc_w_4_000_s_10_000 = 5.77e-12  mcrdlm5p1_cf_w_4_000_s_10_000 = 3.20e-11
+ mcrdlm5p1_ca_w_4_000_s_12_000 = 1.05e-05  mcrdlm5p1_cc_w_4_000_s_12_000 = 3.56e-12  mcrdlm5p1_cf_w_4_000_s_12_000 = 3.40e-11
+ mcrdlm5l1_ca_w_1_600_s_1_600 = 1.13e-05  mcrdlm5l1_cc_w_1_600_s_1_600 = 5.78e-11  mcrdlm5l1_cf_w_1_600_s_1_600 = 9.16e-12
+ mcrdlm5l1_ca_w_1_600_s_1_700 = 1.13e-05  mcrdlm5l1_cc_w_1_600_s_1_700 = 5.49e-11  mcrdlm5l1_cf_w_1_600_s_1_700 = 9.66e-12
+ mcrdlm5l1_ca_w_1_600_s_1_900 = 1.13e-05  mcrdlm5l1_cc_w_1_600_s_1_900 = 4.98e-11  mcrdlm5l1_cf_w_1_600_s_1_900 = 1.06e-11
+ mcrdlm5l1_ca_w_1_600_s_2_000 = 1.13e-05  mcrdlm5l1_cc_w_1_600_s_2_000 = 4.76e-11  mcrdlm5l1_cf_w_1_600_s_2_000 = 1.11e-11
+ mcrdlm5l1_ca_w_1_600_s_2_400 = 1.13e-05  mcrdlm5l1_cc_w_1_600_s_2_400 = 4.03e-11  mcrdlm5l1_cf_w_1_600_s_2_400 = 1.30e-11
+ mcrdlm5l1_ca_w_1_600_s_2_800 = 1.13e-05  mcrdlm5l1_cc_w_1_600_s_2_800 = 3.48e-11  mcrdlm5l1_cf_w_1_600_s_2_800 = 1.48e-11
+ mcrdlm5l1_ca_w_1_600_s_3_200 = 1.13e-05  mcrdlm5l1_cc_w_1_600_s_3_200 = 3.03e-11  mcrdlm5l1_cf_w_1_600_s_3_200 = 1.65e-11
+ mcrdlm5l1_ca_w_1_600_s_4_800 = 1.13e-05  mcrdlm5l1_cc_w_1_600_s_4_800 = 1.86e-11  mcrdlm5l1_cf_w_1_600_s_4_800 = 2.23e-11
+ mcrdlm5l1_ca_w_1_600_s_10_000 = 1.13e-05  mcrdlm5l1_cc_w_1_600_s_10_000 = 4.74e-12  mcrdlm5l1_cf_w_1_600_s_10_000 = 3.25e-11
+ mcrdlm5l1_ca_w_1_600_s_12_000 = 1.13e-05  mcrdlm5l1_cc_w_1_600_s_12_000 = 2.85e-12  mcrdlm5l1_cf_w_1_600_s_12_000 = 3.42e-11
+ mcrdlm5l1_ca_w_4_000_s_1_600 = 1.13e-05  mcrdlm5l1_cc_w_4_000_s_1_600 = 6.15e-11  mcrdlm5l1_cf_w_4_000_s_1_600 = 9.16e-12
+ mcrdlm5l1_ca_w_4_000_s_1_700 = 1.13e-05  mcrdlm5l1_cc_w_4_000_s_1_700 = 5.83e-11  mcrdlm5l1_cf_w_4_000_s_1_700 = 9.66e-12
+ mcrdlm5l1_ca_w_4_000_s_1_900 = 1.13e-05  mcrdlm5l1_cc_w_4_000_s_1_900 = 5.29e-11  mcrdlm5l1_cf_w_4_000_s_1_900 = 1.07e-11
+ mcrdlm5l1_ca_w_4_000_s_2_000 = 1.13e-05  mcrdlm5l1_cc_w_4_000_s_2_000 = 5.06e-11  mcrdlm5l1_cf_w_4_000_s_2_000 = 1.11e-11
+ mcrdlm5l1_ca_w_4_000_s_2_400 = 1.13e-05  mcrdlm5l1_cc_w_4_000_s_2_400 = 4.28e-11  mcrdlm5l1_cf_w_4_000_s_2_400 = 1.30e-11
+ mcrdlm5l1_ca_w_4_000_s_2_800 = 1.13e-05  mcrdlm5l1_cc_w_4_000_s_2_800 = 3.70e-11  mcrdlm5l1_cf_w_4_000_s_2_800 = 1.48e-11
+ mcrdlm5l1_ca_w_4_000_s_3_200 = 1.13e-05  mcrdlm5l1_cc_w_4_000_s_3_200 = 3.22e-11  mcrdlm5l1_cf_w_4_000_s_3_200 = 1.66e-11
+ mcrdlm5l1_ca_w_4_000_s_4_800 = 1.13e-05  mcrdlm5l1_cc_w_4_000_s_4_800 = 1.99e-11  mcrdlm5l1_cf_w_4_000_s_4_800 = 2.25e-11
+ mcrdlm5l1_ca_w_4_000_s_10_000 = 1.13e-05  mcrdlm5l1_cc_w_4_000_s_10_000 = 5.10e-12  mcrdlm5l1_cf_w_4_000_s_10_000 = 3.33e-11
+ mcrdlm5l1_ca_w_4_000_s_12_000 = 1.13e-05  mcrdlm5l1_cc_w_4_000_s_12_000 = 3.11e-12  mcrdlm5l1_cf_w_4_000_s_12_000 = 3.51e-11
+ mcrdlm5m1_ca_w_1_600_s_1_600 = 1.26e-05  mcrdlm5m1_cc_w_1_600_s_1_600 = 5.65e-11  mcrdlm5m1_cf_w_1_600_s_1_600 = 1.02e-11
+ mcrdlm5m1_ca_w_1_600_s_1_700 = 1.26e-05  mcrdlm5m1_cc_w_1_600_s_1_700 = 5.35e-11  mcrdlm5m1_cf_w_1_600_s_1_700 = 1.07e-11
+ mcrdlm5m1_ca_w_1_600_s_1_900 = 1.26e-05  mcrdlm5m1_cc_w_1_600_s_1_900 = 4.85e-11  mcrdlm5m1_cf_w_1_600_s_1_900 = 1.18e-11
+ mcrdlm5m1_ca_w_1_600_s_2_000 = 1.26e-05  mcrdlm5m1_cc_w_1_600_s_2_000 = 4.62e-11  mcrdlm5m1_cf_w_1_600_s_2_000 = 1.23e-11
+ mcrdlm5m1_ca_w_1_600_s_2_400 = 1.26e-05  mcrdlm5m1_cc_w_1_600_s_2_400 = 3.90e-11  mcrdlm5m1_cf_w_1_600_s_2_400 = 1.44e-11
+ mcrdlm5m1_ca_w_1_600_s_2_800 = 1.26e-05  mcrdlm5m1_cc_w_1_600_s_2_800 = 3.33e-11  mcrdlm5m1_cf_w_1_600_s_2_800 = 1.63e-11
+ mcrdlm5m1_ca_w_1_600_s_3_200 = 1.26e-05  mcrdlm5m1_cc_w_1_600_s_3_200 = 2.88e-11  mcrdlm5m1_cf_w_1_600_s_3_200 = 1.81e-11
+ mcrdlm5m1_ca_w_1_600_s_4_800 = 1.26e-05  mcrdlm5m1_cc_w_1_600_s_4_800 = 1.73e-11  mcrdlm5m1_cf_w_1_600_s_4_800 = 2.43e-11
+ mcrdlm5m1_ca_w_1_600_s_10_000 = 1.26e-05  mcrdlm5m1_cc_w_1_600_s_10_000 = 3.98e-12  mcrdlm5m1_cf_w_1_600_s_10_000 = 3.44e-11
+ mcrdlm5m1_ca_w_1_600_s_12_000 = 1.26e-05  mcrdlm5m1_cc_w_1_600_s_12_000 = 2.30e-12  mcrdlm5m1_cf_w_1_600_s_12_000 = 3.59e-11
+ mcrdlm5m1_ca_w_4_000_s_1_600 = 1.26e-05  mcrdlm5m1_cc_w_4_000_s_1_600 = 5.98e-11  mcrdlm5m1_cf_w_4_000_s_1_600 = 1.02e-11
+ mcrdlm5m1_ca_w_4_000_s_1_700 = 1.26e-05  mcrdlm5m1_cc_w_4_000_s_1_700 = 5.66e-11  mcrdlm5m1_cf_w_4_000_s_1_700 = 1.07e-11
+ mcrdlm5m1_ca_w_4_000_s_1_900 = 1.26e-05  mcrdlm5m1_cc_w_4_000_s_1_900 = 5.12e-11  mcrdlm5m1_cf_w_4_000_s_1_900 = 1.18e-11
+ mcrdlm5m1_ca_w_4_000_s_2_000 = 1.26e-05  mcrdlm5m1_cc_w_4_000_s_2_000 = 4.88e-11  mcrdlm5m1_cf_w_4_000_s_2_000 = 1.23e-11
+ mcrdlm5m1_ca_w_4_000_s_2_400 = 1.26e-05  mcrdlm5m1_cc_w_4_000_s_2_400 = 4.11e-11  mcrdlm5m1_cf_w_4_000_s_2_400 = 1.44e-11
+ mcrdlm5m1_ca_w_4_000_s_2_800 = 1.26e-05  mcrdlm5m1_cc_w_4_000_s_2_800 = 3.53e-11  mcrdlm5m1_cf_w_4_000_s_2_800 = 1.64e-11
+ mcrdlm5m1_ca_w_4_000_s_3_200 = 1.26e-05  mcrdlm5m1_cc_w_4_000_s_3_200 = 3.05e-11  mcrdlm5m1_cf_w_4_000_s_3_200 = 1.82e-11
+ mcrdlm5m1_ca_w_4_000_s_4_800 = 1.26e-05  mcrdlm5m1_cc_w_4_000_s_4_800 = 1.83e-11  mcrdlm5m1_cf_w_4_000_s_4_800 = 2.45e-11
+ mcrdlm5m1_ca_w_4_000_s_10_000 = 1.26e-05  mcrdlm5m1_cc_w_4_000_s_10_000 = 4.29e-12  mcrdlm5m1_cf_w_4_000_s_10_000 = 3.52e-11
+ mcrdlm5m1_ca_w_4_000_s_12_000 = 1.26e-05  mcrdlm5m1_cc_w_4_000_s_12_000 = 2.48e-12  mcrdlm5m1_cf_w_4_000_s_12_000 = 3.68e-11
+ mcrdlm5m2_ca_w_1_600_s_1_600 = 1.44e-05  mcrdlm5m2_cc_w_1_600_s_1_600 = 5.48e-11  mcrdlm5m2_cf_w_1_600_s_1_600 = 1.15e-11
+ mcrdlm5m2_ca_w_1_600_s_1_700 = 1.44e-05  mcrdlm5m2_cc_w_1_600_s_1_700 = 5.18e-11  mcrdlm5m2_cf_w_1_600_s_1_700 = 1.22e-11
+ mcrdlm5m2_ca_w_1_600_s_1_900 = 1.44e-05  mcrdlm5m2_cc_w_1_600_s_1_900 = 4.68e-11  mcrdlm5m2_cf_w_1_600_s_1_900 = 1.34e-11
+ mcrdlm5m2_ca_w_1_600_s_2_000 = 1.44e-05  mcrdlm5m2_cc_w_1_600_s_2_000 = 4.45e-11  mcrdlm5m2_cf_w_1_600_s_2_000 = 1.40e-11
+ mcrdlm5m2_ca_w_1_600_s_2_400 = 1.44e-05  mcrdlm5m2_cc_w_1_600_s_2_400 = 3.72e-11  mcrdlm5m2_cf_w_1_600_s_2_400 = 1.62e-11
+ mcrdlm5m2_ca_w_1_600_s_2_800 = 1.44e-05  mcrdlm5m2_cc_w_1_600_s_2_800 = 3.16e-11  mcrdlm5m2_cf_w_1_600_s_2_800 = 1.84e-11
+ mcrdlm5m2_ca_w_1_600_s_3_200 = 1.44e-05  mcrdlm5m2_cc_w_1_600_s_3_200 = 2.70e-11  mcrdlm5m2_cf_w_1_600_s_3_200 = 2.04e-11
+ mcrdlm5m2_ca_w_1_600_s_4_800 = 1.44e-05  mcrdlm5m2_cc_w_1_600_s_4_800 = 1.56e-11  mcrdlm5m2_cf_w_1_600_s_4_800 = 2.69e-11
+ mcrdlm5m2_ca_w_1_600_s_10_000 = 1.44e-05  mcrdlm5m2_cc_w_1_600_s_10_000 = 3.18e-12  mcrdlm5m2_cf_w_1_600_s_10_000 = 3.68e-11
+ mcrdlm5m2_ca_w_1_600_s_12_000 = 1.44e-05  mcrdlm5m2_cc_w_1_600_s_12_000 = 1.75e-12  mcrdlm5m2_cf_w_1_600_s_12_000 = 3.81e-11
+ mcrdlm5m2_ca_w_4_000_s_1_600 = 1.44e-05  mcrdlm5m2_cc_w_4_000_s_1_600 = 5.78e-11  mcrdlm5m2_cf_w_4_000_s_1_600 = 1.15e-11
+ mcrdlm5m2_ca_w_4_000_s_1_700 = 1.44e-05  mcrdlm5m2_cc_w_4_000_s_1_700 = 5.46e-11  mcrdlm5m2_cf_w_4_000_s_1_700 = 1.22e-11
+ mcrdlm5m2_ca_w_4_000_s_1_900 = 1.44e-05  mcrdlm5m2_cc_w_4_000_s_1_900 = 4.92e-11  mcrdlm5m2_cf_w_4_000_s_1_900 = 1.34e-11
+ mcrdlm5m2_ca_w_4_000_s_2_000 = 1.44e-05  mcrdlm5m2_cc_w_4_000_s_2_000 = 4.68e-11  mcrdlm5m2_cf_w_4_000_s_2_000 = 1.40e-11
+ mcrdlm5m2_ca_w_4_000_s_2_400 = 1.44e-05  mcrdlm5m2_cc_w_4_000_s_2_400 = 3.91e-11  mcrdlm5m2_cf_w_4_000_s_2_400 = 1.63e-11
+ mcrdlm5m2_ca_w_4_000_s_2_800 = 1.44e-05  mcrdlm5m2_cc_w_4_000_s_2_800 = 3.32e-11  mcrdlm5m2_cf_w_4_000_s_2_800 = 1.84e-11
+ mcrdlm5m2_ca_w_4_000_s_3_200 = 1.44e-05  mcrdlm5m2_cc_w_4_000_s_3_200 = 2.85e-11  mcrdlm5m2_cf_w_4_000_s_3_200 = 2.04e-11
+ mcrdlm5m2_ca_w_4_000_s_4_800 = 1.44e-05  mcrdlm5m2_cc_w_4_000_s_4_800 = 1.66e-11  mcrdlm5m2_cf_w_4_000_s_4_800 = 2.72e-11
+ mcrdlm5m2_ca_w_4_000_s_10_000 = 1.44e-05  mcrdlm5m2_cc_w_4_000_s_10_000 = 3.46e-12  mcrdlm5m2_cf_w_4_000_s_10_000 = 3.75e-11
+ mcrdlm5m2_ca_w_4_000_s_12_000 = 1.44e-05  mcrdlm5m2_cc_w_4_000_s_12_000 = 1.93e-12  mcrdlm5m2_cf_w_4_000_s_12_000 = 3.90e-11
+ mcrdlm5m3_ca_w_1_600_s_1_600 = 2.10e-05  mcrdlm5m3_cc_w_1_600_s_1_600 = 5.01e-11  mcrdlm5m3_cf_w_1_600_s_1_600 = 1.62e-11
+ mcrdlm5m3_ca_w_1_600_s_1_700 = 2.10e-05  mcrdlm5m3_cc_w_1_600_s_1_700 = 4.71e-11  mcrdlm5m3_cf_w_1_600_s_1_700 = 1.70e-11
+ mcrdlm5m3_ca_w_1_600_s_1_900 = 2.10e-05  mcrdlm5m3_cc_w_1_600_s_1_900 = 4.19e-11  mcrdlm5m3_cf_w_1_600_s_1_900 = 1.87e-11
+ mcrdlm5m3_ca_w_1_600_s_2_000 = 2.10e-05  mcrdlm5m3_cc_w_1_600_s_2_000 = 3.97e-11  mcrdlm5m3_cf_w_1_600_s_2_000 = 1.94e-11
+ mcrdlm5m3_ca_w_1_600_s_2_400 = 2.10e-05  mcrdlm5m3_cc_w_1_600_s_2_400 = 3.24e-11  mcrdlm5m3_cf_w_1_600_s_2_400 = 2.23e-11
+ mcrdlm5m3_ca_w_1_600_s_2_800 = 2.10e-05  mcrdlm5m3_cc_w_1_600_s_2_800 = 2.68e-11  mcrdlm5m3_cf_w_1_600_s_2_800 = 2.50e-11
+ mcrdlm5m3_ca_w_1_600_s_3_200 = 2.10e-05  mcrdlm5m3_cc_w_1_600_s_3_200 = 2.25e-11  mcrdlm5m3_cf_w_1_600_s_3_200 = 2.74e-11
+ mcrdlm5m3_ca_w_1_600_s_4_800 = 2.10e-05  mcrdlm5m3_cc_w_1_600_s_4_800 = 1.17e-11  mcrdlm5m3_cf_w_1_600_s_4_800 = 3.47e-11
+ mcrdlm5m3_ca_w_1_600_s_10_000 = 2.10e-05  mcrdlm5m3_cc_w_1_600_s_10_000 = 1.81e-12  mcrdlm5m3_cf_w_1_600_s_10_000 = 4.33e-11
+ mcrdlm5m3_ca_w_1_600_s_12_000 = 2.10e-05  mcrdlm5m3_cc_w_1_600_s_12_000 = 9.00e-13  mcrdlm5m3_cf_w_1_600_s_12_000 = 4.42e-11
+ mcrdlm5m3_ca_w_4_000_s_1_600 = 2.10e-05  mcrdlm5m3_cc_w_4_000_s_1_600 = 5.23e-11  mcrdlm5m3_cf_w_4_000_s_1_600 = 1.62e-11
+ mcrdlm5m3_ca_w_4_000_s_1_700 = 2.10e-05  mcrdlm5m3_cc_w_4_000_s_1_700 = 4.92e-11  mcrdlm5m3_cf_w_4_000_s_1_700 = 1.70e-11
+ mcrdlm5m3_ca_w_4_000_s_1_900 = 2.10e-05  mcrdlm5m3_cc_w_4_000_s_1_900 = 4.39e-11  mcrdlm5m3_cf_w_4_000_s_1_900 = 1.87e-11
+ mcrdlm5m3_ca_w_4_000_s_2_000 = 2.10e-05  mcrdlm5m3_cc_w_4_000_s_2_000 = 4.15e-11  mcrdlm5m3_cf_w_4_000_s_2_000 = 1.95e-11
+ mcrdlm5m3_ca_w_4_000_s_2_400 = 2.10e-05  mcrdlm5m3_cc_w_4_000_s_2_400 = 3.39e-11  mcrdlm5m3_cf_w_4_000_s_2_400 = 2.24e-11
+ mcrdlm5m3_ca_w_4_000_s_2_800 = 2.10e-05  mcrdlm5m3_cc_w_4_000_s_2_800 = 2.82e-11  mcrdlm5m3_cf_w_4_000_s_2_800 = 2.51e-11
+ mcrdlm5m3_ca_w_4_000_s_3_200 = 2.10e-05  mcrdlm5m3_cc_w_4_000_s_3_200 = 2.37e-11  mcrdlm5m3_cf_w_4_000_s_3_200 = 2.75e-11
+ mcrdlm5m3_ca_w_4_000_s_4_800 = 2.10e-05  mcrdlm5m3_cc_w_4_000_s_4_800 = 1.26e-11  mcrdlm5m3_cf_w_4_000_s_4_800 = 3.50e-11
+ mcrdlm5m3_ca_w_4_000_s_10_000 = 2.10e-05  mcrdlm5m3_cc_w_4_000_s_10_000 = 1.98e-12  mcrdlm5m3_cf_w_4_000_s_10_000 = 4.40e-11
+ mcrdlm5m3_ca_w_4_000_s_12_000 = 2.10e-05  mcrdlm5m3_cc_w_4_000_s_12_000 = 9.85e-13  mcrdlm5m3_cf_w_4_000_s_12_000 = 4.50e-11
+ mcrdlm5m4_ca_w_1_600_s_1_600 = 5.30e-05  mcrdlm5m4_cc_w_1_600_s_1_600 = 3.92e-11  mcrdlm5m4_cf_w_1_600_s_1_600 = 3.42e-11
+ mcrdlm5m4_ca_w_1_600_s_1_700 = 5.30e-05  mcrdlm5m4_cc_w_1_600_s_1_700 = 3.63e-11  mcrdlm5m4_cf_w_1_600_s_1_700 = 3.56e-11
+ mcrdlm5m4_ca_w_1_600_s_1_900 = 5.30e-05  mcrdlm5m4_cc_w_1_600_s_1_900 = 3.14e-11  mcrdlm5m4_cf_w_1_600_s_1_900 = 3.80e-11
+ mcrdlm5m4_ca_w_1_600_s_2_000 = 5.30e-05  mcrdlm5m4_cc_w_1_600_s_2_000 = 2.93e-11  mcrdlm5m4_cf_w_1_600_s_2_000 = 3.92e-11
+ mcrdlm5m4_ca_w_1_600_s_2_400 = 5.30e-05  mcrdlm5m4_cc_w_1_600_s_2_400 = 2.26e-11  mcrdlm5m4_cf_w_1_600_s_2_400 = 4.34e-11
+ mcrdlm5m4_ca_w_1_600_s_2_800 = 5.30e-05  mcrdlm5m4_cc_w_1_600_s_2_800 = 1.78e-11  mcrdlm5m4_cf_w_1_600_s_2_800 = 4.67e-11
+ mcrdlm5m4_ca_w_1_600_s_3_200 = 5.30e-05  mcrdlm5m4_cc_w_1_600_s_3_200 = 1.42e-11  mcrdlm5m4_cf_w_1_600_s_3_200 = 4.94e-11
+ mcrdlm5m4_ca_w_1_600_s_4_800 = 5.30e-05  mcrdlm5m4_cc_w_1_600_s_4_800 = 6.24e-12  mcrdlm5m4_cf_w_1_600_s_4_800 = 5.61e-11
+ mcrdlm5m4_ca_w_1_600_s_10_000 = 5.30e-05  mcrdlm5m4_cc_w_1_600_s_10_000 = 6.60e-13  mcrdlm5m4_cf_w_1_600_s_10_000 = 6.13e-11
+ mcrdlm5m4_ca_w_1_600_s_12_000 = 5.30e-05  mcrdlm5m4_cc_w_1_600_s_12_000 = 2.95e-13  mcrdlm5m4_cf_w_1_600_s_12_000 = 6.17e-11
+ mcrdlm5m4_ca_w_4_000_s_1_600 = 5.30e-05  mcrdlm5m4_cc_w_4_000_s_1_600 = 4.13e-11  mcrdlm5m4_cf_w_4_000_s_1_600 = 3.43e-11
+ mcrdlm5m4_ca_w_4_000_s_1_700 = 5.30e-05  mcrdlm5m4_cc_w_4_000_s_1_700 = 3.82e-11  mcrdlm5m4_cf_w_4_000_s_1_700 = 3.56e-11
+ mcrdlm5m4_ca_w_4_000_s_1_900 = 5.30e-05  mcrdlm5m4_cc_w_4_000_s_1_900 = 3.33e-11  mcrdlm5m4_cf_w_4_000_s_1_900 = 3.81e-11
+ mcrdlm5m4_ca_w_4_000_s_2_000 = 5.30e-05  mcrdlm5m4_cc_w_4_000_s_2_000 = 3.12e-11  mcrdlm5m4_cf_w_4_000_s_2_000 = 3.93e-11
+ mcrdlm5m4_ca_w_4_000_s_2_400 = 5.30e-05  mcrdlm5m4_cc_w_4_000_s_2_400 = 2.41e-11  mcrdlm5m4_cf_w_4_000_s_2_400 = 4.34e-11
+ mcrdlm5m4_ca_w_4_000_s_2_800 = 5.30e-05  mcrdlm5m4_cc_w_4_000_s_2_800 = 1.91e-11  mcrdlm5m4_cf_w_4_000_s_2_800 = 4.68e-11
+ mcrdlm5m4_ca_w_4_000_s_3_200 = 5.30e-05  mcrdlm5m4_cc_w_4_000_s_3_200 = 1.53e-11  mcrdlm5m4_cf_w_4_000_s_3_200 = 4.96e-11
+ mcrdlm5m4_ca_w_4_000_s_4_800 = 5.30e-05  mcrdlm5m4_cc_w_4_000_s_4_800 = 6.98e-12  mcrdlm5m4_cf_w_4_000_s_4_800 = 5.65e-11
+ mcrdlm5m4_ca_w_4_000_s_10_000 = 5.30e-05  mcrdlm5m4_cc_w_4_000_s_10_000 = 8.05e-13  mcrdlm5m4_cf_w_4_000_s_10_000 = 6.24e-11
+ mcrdlm5m4_ca_w_4_000_s_12_000 = 5.30e-05  mcrdlm5m4_cc_w_4_000_s_12_000 = 3.75e-13  mcrdlm5m4_cf_w_4_000_s_12_000 = 6.28e-11
+ cp1f = 8.04e-05  cp1fsw = 7.43e-11
+ cl1f = 2.93e-05  cl1fsw = 6.80e-11
+ cl1d = 4.53e-05  cl1dsw = 6.75e-11
+ cl1p1 = 6.45e-05  cl1p1sw = 6.70e-11
+ cm1f = 2.02e-05  cm1fsw = 8.97e-11
+ cm1d = 2.67e-05  cm1dsw = 8.96e-11
+ cm1p1 = 3.23e-05  cm1p1sw = 8.92e-11
+ cm1l1 = 7.72e-05  cm1l1sw = 8.81e-11
+ cm2f = 1.40e-05  cm2fsw = 8.98e-11
+ cm2d = 1.68e-05  cm2dsw = 8.98e-11
+ cm2p1 = 1.89e-05  cm2p1sw = 8.95e-11
+ cm2l1 = 2.86e-05  cm2l1sw = 8.92e-11
+ cm2m1 = 8.04e-05  cm2m1sw = 8.78e-11
+ cm3f = 1.02e-05  cm3fsw = 9.37e-11
+ cm3d = 1.17e-05  cm3dsw = 9.35e-11
+ cm3p1 = 1.26e-05  cm3p1sw = 9.35e-11
+ cm3l1 = 1.63e-05  cm3l1sw = 9.31e-11
+ cm3m1 = 2.58e-05  cm3m1sw = 9.25e-11
+ cm3m2 = 5.95e-05  cm3m2sw = 9.12e-11
+ cm4f = 7.28e-06  cm4fsw = 9.41e-11
+ cm4d = 7.98e-06  cm4dsw = 9.40e-11
+ cm4p1 = 8.42e-06  cm4p1sw = 9.40e-11
+ cm4l1 = 9.92e-06  cm4l1sw = 9.38e-11
+ cm4m1 = 1.28e-05  cm4m1sw = 9.36e-11
+ cm4m2 = 1.78e-05  cm4m2sw = 9.32e-11
+ cm4m3 = 5.76e-05  cm4m3sw = 9.14e-11
+ cm5f = 5.56e-06  cm5fsw = 6.93e-11
+ cm5d = 5.96e-06  cm5dsw = 6.91e-11
+ cm5p1 = 6.20e-06  cm5p1sw = 6.92e-11
+ cm5l1 = 6.97e-06  cm5l1sw = 6.90e-11
+ cm5m1 = 8.26e-06  cm5m1sw = 6.86e-11
+ cm5m2 = 1.01e-05  cm5m2sw = 6.84e-11
+ cm5m3 = 1.67e-05  cm5m3sw = 6.82e-11
+ cm5m4 = 4.87e-05  cm5m4sw = 7.53e-11
+ crdlf = 2.15e-06  crdlfsw = 4.71e-11
+ crdld = 2.21e-06  crdldsw = 4.71e-11
+ crdlp1 = 2.24e-06  crdlp1sw = 4.70e-11
+ crdll1 = 2.33e-06  crdll1sw = 4.69e-11
+ crdlm1 = 2.46e-06  crdlm1sw = 4.68e-11
+ crdlm2 = 2.60e-06  crdlm2sw = 4.67e-11
+ crdlm3 = 2.90e-06  crdlm3sw = 4.65e-11
+ crdlm4 = 3.28e-06  crdlm4sw = 4.64e-11
+ crdlm5 = 4.28e-06  crdlm5sw = 4.65e-11
+ cl1p1f = 1.45e-04  cl1p1fsw = 7.25e-11
+ cm1p1f = 1.13e-04  cm1p1fsw = 7.33e-11
+ cm2p1f = 9.94e-05  cm2p1fsw = 7.38e-11
+ cm3p1f = 9.31e-05  cm3p1fsw = 7.40e-11
+ cm4p1f = 8.89e-05  cm4p1fsw = 7.42e-11
+ cm5p1f = 8.66e-05  cm5p1fsw = 7.42e-11
+ crdlp1f = 8.27e-05  crdlp1fsw = 7.43e-11
+ cm1l1f = 1.07e-04  cm1l1fsw = 6.58e-11
+ cm1l1d = 1.23e-04  cm1l1dsw = 6.52e-11
+ cm1l1p1 = 1.42e-04  cm1l1p1sw = 6.47e-11
+ cm2l1f = 5.80e-05  cm2l1fsw = 6.71e-11
+ cm2l1d = 7.39e-05  cm2l1dsw = 6.66e-11
+ cm2l1p1 = 9.32e-05  cm2l1p1sw = 6.61e-11
+ cm3l1f = 4.57e-05  cm3l1fsw = 6.76e-11
+ cm3l1d = 6.16e-05  cm3l1dsw = 6.71e-11
+ cm3l1p1 = 8.09e-05  cm3l1p1sw = 6.66e-11
+ cm4l1f = 3.93e-05  cm4l1fsw = 6.79e-11
+ cm4l1d = 5.52e-05  cm4l1dsw = 6.73e-11
+ cm4l1p1 = 7.44e-05  cm4l1p1sw = 6.68e-11
+ cm5l1f = 3.63e-05  cm5l1fsw = 6.80e-11
+ cm5l1d = 5.22e-05  cm5l1dsw = 6.73e-11
+ cm5l1p1 = 7.15e-05  cm5l1p1sw = 6.69e-11
+ crdll1f = 3.17e-05  crdll1fsw = 6.80e-11
+ crdll1d = 4.76e-05  crdll1dsw = 6.74e-11
+ crdll1p1 = 6.68e-05  crdll1p1sw = 6.70e-11
+ cm2m1f = 1.01e-04  cm2m1fsw = 8.77e-11
+ cm2m1d = 1.07e-04  cm2m1dsw = 8.75e-11
+ cm2m1p1 = 1.13e-04  cm2m1p1sw = 8.73e-11
+ cm2m1l1 = 1.58e-04  cm2m1l1sw = 8.58e-11
+ cm3m1f = 4.60e-05  cm3m1fsw = 8.87e-11
+ cm3m1d = 5.25e-05  cm3m1dsw = 8.81e-11
+ cm3m1p1 = 5.81e-05  cm3m1p1sw = 8.80e-11
+ cm3m1l1 = 1.03e-04  cm3m1l1sw = 8.73e-11
+ cm4m1f = 3.30e-05  cm4m1fsw = 8.93e-11
+ cm4m1d = 3.94e-05  cm4m1dsw = 8.91e-11
+ cm4m1p1 = 4.51e-05  cm4m1p1sw = 8.91e-11
+ cm4m1l1 = 9.00e-05  cm4m1l1sw = 8.79e-11
+ cm5m1f = 2.85e-05  cm5m1fsw = 8.94e-11
+ cm5m1d = 3.49e-05  cm5m1dsw = 8.92e-11
+ cm5m1p1 = 4.06e-05  cm5m1p1sw = 8.91e-11
+ cm5m1l1 = 8.55e-05  cm5m1l1sw = 8.81e-11
+ crdlm1f = 2.27e-05  crdlm1fsw = 8.98e-11
+ crdlm1d = 2.91e-05  crdlm1dsw = 8.96e-11
+ crdlm1p1 = 3.48e-05  crdlm1p1sw = 8.93e-11
+ crdlm1l1 = 7.97e-05  crdlm1l1sw = 8.82e-11
+ cm3m2f = 7.34e-05  cm3m2fsw = 8.83e-11
+ cm3m2d = 7.63e-05  cm3m2dsw = 8.83e-11
+ cm3m2p1 = 7.84e-05  cm3m2p1sw = 8.82e-11
+ cm3m2l1 = 8.81e-05  cm3m2l1sw = 8.79e-11
+ cm3m2m1 = 1.40e-04  cm3m2m1sw = 8.59e-11
+ cm4m2f = 3.17e-05  cm4m2fsw = 8.96e-11
+ cm4m2d = 3.46e-05  cm4m2dsw = 8.91e-11
+ cm4m2p1 = 3.67e-05  cm4m2p1sw = 8.93e-11
+ cm4m2l1 = 4.64e-05  cm4m2l1sw = 8.87e-11
+ cm4m2m1 = 9.81e-05  cm4m2m1sw = 8.77e-11
+ cm5m2f = 2.41e-05  cm5m2fsw = 9.01e-11
+ cm5m2d = 2.69e-05  cm5m2dsw = 9.00e-11
+ cm5m2p1 = 2.90e-05  cm5m2p1sw = 9.00e-11
+ cm5m2l1 = 3.87e-05  cm5m2l1sw = 8.90e-11
+ cm5m2m1 = 9.05e-05  cm5m2m1sw = 8.80e-11
+ crdlm2f = 1.66e-05  crdlm2fsw = 8.99e-11
+ crdlm2d = 1.94e-05  crdlm2dsw = 8.98e-11
+ crdlm2p1 = 2.15e-05  crdlm2p1sw = 8.96e-11
+ crdlm2l1 = 3.12e-05  crdlm2l1sw = 8.93e-11
+ crdlm2m1 = 8.30e-05  crdlm2m1sw = 8.83e-11
+ cm4m3f = 6.78e-05  cm4m3fsw = 9.08e-11
+ cm4m3d = 6.92e-05  cm4m3dsw = 9.06e-11
+ cm4m3p1 = 7.02e-05  cm4m3p1sw = 9.03e-11
+ cm4m3l1 = 7.39e-05  cm4m3l1sw = 9.03e-11
+ cm4m3m1 = 8.33e-05  cm4m3m1sw = 8.96e-11
+ cm4m3m2 = 1.17e-04  cm4m3m2sw = 8.83e-11
+ cm5m3f = 2.69e-05  cm5m3fsw = 9.23e-11
+ cm5m3d = 2.83e-05  cm5m3dsw = 9.21e-11
+ cm5m3p1 = 2.93e-05  cm5m3p1sw = 9.21e-11
+ cm5m3l1 = 3.30e-05  cm5m3l1sw = 9.17e-11
+ cm5m3m1 = 4.24e-05  cm5m3m1sw = 9.11e-11
+ cm5m3m2 = 7.61e-05  cm5m3m2sw = 9.01e-11
+ crdlm3f = 1.31e-05  crdlm3fsw = 9.37e-11
+ crdlm3d = 1.45e-05  crdlm3dsw = 9.37e-11
+ crdlm3p1 = 1.55e-05  crdlm3p1sw = 9.36e-11
+ crdlm3l1 = 1.92e-05  crdlm3l1sw = 9.32e-11
+ crdlm3m1 = 2.87e-05  crdlm3m1sw = 9.24e-11
+ crdlm3m2 = 6.23e-05  crdlm3m2sw = 9.14e-11
+ cm5m4f = 5.59e-05  cm5m4fsw = 9.12e-11
+ cm5m4d = 5.66e-05  cm5m4dsw = 9.11e-11
+ cm5m4p1 = 5.71e-05  cm5m4p1sw = 9.09e-11
+ cm5m4l1 = 5.86e-05  cm5m4l1sw = 9.07e-11
+ cm5m4m1 = 6.14e-05  cm5m4m1sw = 9.07e-11
+ cm5m4m2 = 6.64e-05  cm5m4m2sw = 9.02e-11
+ cm5m4m3 = 1.06e-04  cm5m4m3sw = 8.86e-11
+ crdlm4f = 1.06e-05  crdlm4fsw = 9.42e-11
+ crdlm4d = 1.12e-05  crdlm4dsw = 9.42e-11
+ crdlm4p1 = 1.17e-05  crdlm4p1sw = 9.41e-11
+ crdlm4l1 = 1.32e-05  crdlm4l1sw = 9.40e-11
+ crdlm4m1 = 1.60e-05  crdlm4m1sw = 9.36e-11
+ crdlm4m2 = 2.10e-05  crdlm4m2sw = 9.30e-11
+ crdlm4m3 = 6.09e-05  crdlm4m3sw = 9.14e-11
+ crdlm5f = 9.86e-06  crdlm5fsw = 6.75e-11
+ crdlm5d = 1.03e-05  crdlm5dsw = 6.73e-11
+ crdlm5p1 = 1.05e-05  crdlm5p1sw = 6.72e-11
+ crdlm5l1 = 1.13e-05  crdlm5l1sw = 6.70e-11
+ crdlm5m1 = 1.26e-05  crdlm5m1sw = 6.67e-11
+ crdlm5m2 = 1.44e-05  crdlm5m2sw = 6.64e-11
+ crdlm5m3 = 2.10e-05  crdlm5m3sw = 6.63e-11
+ crdlm5m4 = 5.30e-05  crdlm5m4sw = 7.34e-11
