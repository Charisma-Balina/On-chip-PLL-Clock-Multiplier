* SKY130 Spice File.
.param
+ tol_nfom=-0.069u
+ tol_pfom=-0.060u
+ tol_nw = -0.069u
+ tol_poly = -0.041u
+ tol_li = -0.020u
+ tol_m1 = -0.025u
+ tol_m2 = -0.025u
+ tol_m3 = -0.065u
+ tol_m4 = -0.065u
+ tol_m5 = -0.17u
+ tol_rdl = -1.0u
.param
+ rcn=345
+ rcp=870
+ rdn=132
+ rdp=228
+ rdn_hv=126
+ rdp_hv=222
+ rp1=55.80
+ rnw=2160
+ rl1=14.8
+ rm1=0.145
+ rm2=0.145
+ rm3=0.056
+ rm4=0.056
+ rm5=0.0358
+ rrdl=0.0067
+ rcp1=243.28
+ rcl1=22.6
+ rcvia=15
+ rcvia2=8
+ rcvia3=8
+ rcvia4=0.891
+ rcrdlcon=0.0077
+ rspwres=4829
* P+ Poly Preres Parameters
.param
+ crpf_precision=  8.09e-5   $ Units: farad/meter^2
+ crpfsw_precision_1_1 = 4.51e-11 $ Units: farad/meter
+ crpfsw_precision_2_1 = 4.86e-11 $ Units: farad/meter
+ crpfsw_precision_4_1 = 5.28e-11 $ Units: farad/meter
+ crpfsw_precision_8_2 = 5.79e-11 $ Units: farad/meter
+ crpfsw_precision_16_2 = 6.36e-11 $ Units: farad/meter
.include "../sky130_fd_pr__model__r+c.model.spice"
.include "../parameters/fast.spice"
