magic
tech sky130A
timestamp 1605977318
<< nwell >>
rect 374 344 902 640
rect 48 235 902 344
<< nmos >>
rect 48 462 63 546
rect 119 408 227 423
rect 138 144 153 186
rect 238 144 253 186
rect 338 144 353 186
rect 438 144 453 186
rect 538 144 553 186
rect 638 144 653 186
rect 738 66 753 186
rect 840 133 855 187
<< pmos >>
rect 570 461 585 545
rect 688 527 703 569
rect 393 403 501 418
rect 138 253 153 295
rect 238 253 253 295
rect 338 253 353 295
rect 438 253 453 295
rect 538 253 553 295
rect 638 253 653 295
rect 738 253 753 493
rect 840 253 855 361
<< ndiff >>
rect 19 524 48 546
rect 19 506 25 524
rect 42 506 48 524
rect 19 488 48 506
rect 19 470 25 488
rect 42 470 48 488
rect 19 462 48 470
rect 63 523 92 546
rect 63 506 69 523
rect 86 506 92 523
rect 63 488 92 506
rect 63 470 69 488
rect 86 470 92 488
rect 63 462 92 470
rect 119 446 227 452
rect 119 429 127 446
rect 144 429 161 446
rect 178 429 195 446
rect 212 429 227 446
rect 119 423 227 429
rect 119 402 227 408
rect 119 385 123 402
rect 140 385 157 402
rect 174 385 191 402
rect 208 385 227 402
rect 119 379 227 385
rect 109 173 138 186
rect 109 156 115 173
rect 132 156 138 173
rect 109 144 138 156
rect 153 173 182 186
rect 153 156 159 173
rect 176 156 182 173
rect 153 144 182 156
rect 209 173 238 186
rect 209 156 215 173
rect 232 156 238 173
rect 209 144 238 156
rect 253 173 282 186
rect 253 156 259 173
rect 276 156 282 173
rect 253 144 282 156
rect 309 173 338 186
rect 309 156 315 173
rect 332 156 338 173
rect 309 144 338 156
rect 353 173 382 186
rect 353 156 359 173
rect 376 156 382 173
rect 353 144 382 156
rect 409 173 438 186
rect 409 156 415 173
rect 432 156 438 173
rect 409 144 438 156
rect 453 173 482 186
rect 453 156 459 173
rect 476 156 482 173
rect 453 144 482 156
rect 509 173 538 186
rect 509 156 515 173
rect 532 156 538 173
rect 509 144 538 156
rect 553 173 582 186
rect 553 156 559 173
rect 576 156 582 173
rect 553 144 582 156
rect 609 173 638 186
rect 609 156 615 173
rect 632 156 638 173
rect 609 144 638 156
rect 653 173 682 186
rect 653 156 659 173
rect 676 156 682 173
rect 653 144 682 156
rect 709 173 738 186
rect 709 156 715 173
rect 732 156 738 173
rect 709 139 738 156
rect 709 122 715 139
rect 732 122 738 139
rect 709 105 738 122
rect 709 88 715 105
rect 732 88 738 105
rect 709 66 738 88
rect 753 173 782 186
rect 753 156 759 173
rect 776 156 782 173
rect 753 139 782 156
rect 753 122 759 139
rect 776 122 782 139
rect 811 167 840 187
rect 811 150 817 167
rect 834 150 840 167
rect 811 133 840 150
rect 855 167 884 187
rect 855 150 861 167
rect 878 150 884 167
rect 855 133 884 150
rect 753 105 782 122
rect 753 88 759 105
rect 776 88 782 105
rect 753 66 782 88
<< pdiff >>
rect 655 556 688 569
rect 541 537 570 545
rect 541 520 547 537
rect 564 520 570 537
rect 541 503 570 520
rect 541 486 547 503
rect 564 486 570 503
rect 541 461 570 486
rect 585 541 614 545
rect 585 524 591 541
rect 608 524 614 541
rect 655 539 663 556
rect 680 539 688 556
rect 655 527 688 539
rect 703 556 736 569
rect 703 539 711 556
rect 728 539 736 556
rect 703 527 736 539
rect 585 507 614 524
rect 585 490 591 507
rect 608 490 614 507
rect 585 461 614 490
rect 393 441 501 447
rect 393 424 401 441
rect 418 424 435 441
rect 452 424 469 441
rect 486 424 501 441
rect 393 418 501 424
rect 709 451 738 493
rect 709 434 715 451
rect 732 434 738 451
rect 709 409 738 434
rect 393 397 501 403
rect 393 380 401 397
rect 418 380 435 397
rect 452 380 469 397
rect 486 380 501 397
rect 393 374 501 380
rect 709 392 715 409
rect 732 392 738 409
rect 709 367 738 392
rect 709 350 715 367
rect 732 350 738 367
rect 709 325 738 350
rect 709 308 715 325
rect 732 308 738 325
rect 109 283 138 295
rect 109 266 115 283
rect 132 266 138 283
rect 109 253 138 266
rect 153 283 182 295
rect 153 266 159 283
rect 176 266 182 283
rect 153 253 182 266
rect 209 283 238 295
rect 209 266 215 283
rect 232 266 238 283
rect 209 253 238 266
rect 253 283 282 295
rect 253 266 259 283
rect 276 266 282 283
rect 253 253 282 266
rect 309 283 338 295
rect 309 266 315 283
rect 332 266 338 283
rect 309 253 338 266
rect 353 283 382 295
rect 353 266 359 283
rect 376 266 382 283
rect 353 253 382 266
rect 409 283 438 295
rect 409 266 415 283
rect 432 266 438 283
rect 409 253 438 266
rect 453 283 482 295
rect 453 266 459 283
rect 476 266 482 283
rect 453 253 482 266
rect 509 283 538 295
rect 509 266 515 283
rect 532 266 538 283
rect 509 253 538 266
rect 553 283 582 295
rect 553 266 559 283
rect 576 266 582 283
rect 553 253 582 266
rect 609 283 638 295
rect 609 266 615 283
rect 632 266 638 283
rect 609 253 638 266
rect 653 283 682 295
rect 653 266 659 283
rect 676 266 682 283
rect 653 253 682 266
rect 709 283 738 308
rect 709 266 715 283
rect 732 266 738 283
rect 709 253 738 266
rect 753 451 783 493
rect 753 434 759 451
rect 776 434 783 451
rect 753 409 783 434
rect 753 392 759 409
rect 776 392 783 409
rect 753 367 783 392
rect 753 350 759 367
rect 776 350 783 367
rect 753 325 783 350
rect 753 308 759 325
rect 776 308 783 325
rect 753 283 783 308
rect 753 266 759 283
rect 776 266 783 283
rect 753 253 783 266
rect 811 355 840 361
rect 811 337 817 355
rect 834 337 840 355
rect 811 319 840 337
rect 811 301 817 319
rect 834 301 840 319
rect 811 283 840 301
rect 811 266 817 283
rect 834 266 840 283
rect 811 253 840 266
rect 855 348 884 361
rect 855 331 861 348
rect 878 331 884 348
rect 855 313 884 331
rect 855 295 861 313
rect 878 295 884 313
rect 855 277 884 295
rect 855 259 861 277
rect 878 259 884 277
rect 855 253 884 259
<< ndiffc >>
rect 25 506 42 524
rect 25 470 42 488
rect 69 506 86 523
rect 69 470 86 488
rect 127 429 144 446
rect 161 429 178 446
rect 195 429 212 446
rect 123 385 140 402
rect 157 385 174 402
rect 191 385 208 402
rect 115 156 132 173
rect 159 156 176 173
rect 215 156 232 173
rect 259 156 276 173
rect 315 156 332 173
rect 359 156 376 173
rect 415 156 432 173
rect 459 156 476 173
rect 515 156 532 173
rect 559 156 576 173
rect 615 156 632 173
rect 659 156 676 173
rect 715 156 732 173
rect 715 122 732 139
rect 715 88 732 105
rect 759 156 776 173
rect 759 122 776 139
rect 817 150 834 167
rect 861 150 878 167
rect 759 88 776 105
<< pdiffc >>
rect 547 520 564 537
rect 547 486 564 503
rect 591 524 608 541
rect 663 539 680 556
rect 711 539 728 556
rect 591 490 608 507
rect 401 424 418 441
rect 435 424 452 441
rect 469 424 486 441
rect 715 434 732 451
rect 401 380 418 397
rect 435 380 452 397
rect 469 380 486 397
rect 715 392 732 409
rect 715 350 732 367
rect 715 308 732 325
rect 115 266 132 283
rect 159 266 176 283
rect 215 266 232 283
rect 259 266 276 283
rect 315 266 332 283
rect 359 266 376 283
rect 415 266 432 283
rect 459 266 476 283
rect 515 266 532 283
rect 559 266 576 283
rect 615 266 632 283
rect 659 266 676 283
rect 715 266 732 283
rect 759 434 776 451
rect 759 392 776 409
rect 759 350 776 367
rect 759 308 776 325
rect 759 266 776 283
rect 817 337 834 355
rect 817 301 834 319
rect 817 266 834 283
rect 861 331 878 348
rect 861 295 878 313
rect 861 259 878 277
<< psubdiff >>
rect 283 425 295 442
rect 312 425 324 442
rect 283 378 295 395
rect 312 378 324 395
<< nsubdiff >>
rect 408 605 420 622
rect 444 605 456 622
rect 504 605 516 622
rect 540 605 552 622
rect 600 605 612 622
rect 636 605 648 622
rect 696 605 708 622
rect 732 605 744 622
rect 792 605 804 622
rect 828 605 840 622
<< psubdiffcont >>
rect 295 425 312 442
rect 295 378 312 395
<< nsubdiffcont >>
rect 420 605 444 622
rect 516 605 540 622
rect 612 605 636 622
rect 708 605 732 622
rect 804 605 828 622
<< poly >>
rect 48 546 63 559
rect 461 555 585 575
rect 688 569 703 582
rect 461 545 484 555
rect 570 545 585 555
rect 451 534 484 545
rect 451 517 459 534
rect 476 517 484 534
rect 451 512 484 517
rect 48 448 63 462
rect 688 517 703 527
rect 647 502 703 517
rect 647 490 684 502
rect 738 493 753 506
rect 647 473 655 490
rect 673 473 684 490
rect 647 467 684 473
rect 48 447 82 448
rect 47 437 82 447
rect 47 420 55 437
rect 72 423 82 437
rect 72 420 119 423
rect 47 408 119 420
rect 227 408 240 423
rect 570 418 585 461
rect 380 403 393 418
rect 501 403 585 418
rect 138 295 153 308
rect 238 295 253 308
rect 338 295 353 308
rect 438 295 453 308
rect 538 295 553 308
rect 638 295 653 308
rect 840 361 855 374
rect 138 245 153 253
rect 238 245 253 253
rect 338 245 353 253
rect 438 245 453 253
rect 538 245 553 253
rect 638 245 653 253
rect 738 245 753 253
rect 131 235 153 245
rect 231 235 253 245
rect 331 235 353 245
rect 431 235 453 245
rect 531 235 553 245
rect 631 235 653 245
rect 731 235 753 245
rect 109 228 153 235
rect 109 211 117 228
rect 134 211 153 228
rect 109 205 153 211
rect 209 228 253 235
rect 209 211 217 228
rect 234 211 253 228
rect 209 205 253 211
rect 309 228 353 235
rect 309 211 317 228
rect 334 211 353 228
rect 309 205 353 211
rect 409 228 453 235
rect 409 211 417 228
rect 434 211 453 228
rect 409 205 453 211
rect 509 228 553 235
rect 509 211 517 228
rect 534 211 553 228
rect 509 205 553 211
rect 609 228 653 235
rect 609 211 617 228
rect 634 211 653 228
rect 609 205 653 211
rect 709 228 753 235
rect 840 234 855 253
rect 709 211 717 228
rect 734 211 753 228
rect 709 205 753 211
rect 810 228 855 234
rect 810 211 818 228
rect 835 211 855 228
rect 810 205 855 211
rect 131 194 153 205
rect 231 194 253 205
rect 331 194 353 205
rect 431 194 453 205
rect 531 194 553 205
rect 631 194 653 205
rect 731 194 753 205
rect 138 186 153 194
rect 238 186 253 194
rect 338 186 353 194
rect 438 186 453 194
rect 538 186 553 194
rect 638 186 653 194
rect 738 186 753 194
rect 840 187 855 205
rect 138 131 153 144
rect 238 131 253 144
rect 338 131 353 144
rect 438 131 453 144
rect 538 131 553 144
rect 638 131 653 144
rect 840 120 855 133
rect 738 53 753 66
<< polycont >>
rect 459 517 476 534
rect 655 473 673 490
rect 55 420 72 437
rect 117 211 134 228
rect 217 211 234 228
rect 317 211 334 228
rect 417 211 434 228
rect 517 211 534 228
rect 617 211 634 228
rect 717 211 734 228
rect 818 211 835 228
<< locali >>
rect 0 605 12 622
rect 29 605 46 622
rect 63 605 80 622
rect 97 605 114 622
rect 131 605 148 622
rect 165 605 182 622
rect 199 605 216 622
rect 233 605 250 622
rect 267 605 284 622
rect 301 605 318 622
rect 335 605 352 622
rect 369 605 386 622
rect 403 605 420 622
rect 444 605 454 622
rect 471 605 488 622
rect 505 605 516 622
rect 540 605 556 622
rect 573 605 590 622
rect 607 605 612 622
rect 641 605 658 622
rect 675 605 692 622
rect 743 605 760 622
rect 777 605 794 622
rect 845 605 862 622
rect 879 605 902 622
rect 646 556 680 605
rect 25 524 42 546
rect 25 488 42 506
rect 25 462 42 470
rect 69 523 86 546
rect 547 537 564 545
rect 430 534 547 536
rect 430 530 459 534
rect 430 510 436 530
rect 458 517 459 530
rect 476 520 547 534
rect 476 517 564 520
rect 458 510 564 517
rect 69 488 337 506
rect 86 478 337 488
rect 430 503 564 510
rect 430 486 547 503
rect 430 484 564 486
rect 69 462 86 470
rect 139 474 337 478
rect 139 446 209 474
rect 271 449 337 474
rect 547 461 564 484
rect 591 541 611 549
rect 608 512 611 541
rect 646 539 663 556
rect 646 527 680 539
rect 710 556 834 569
rect 710 539 711 556
rect 728 539 834 556
rect 710 527 834 539
rect 591 507 611 512
rect 608 490 611 507
rect 7 437 80 439
rect 7 420 55 437
rect 72 420 80 437
rect 119 429 127 446
rect 144 429 161 446
rect 178 429 195 446
rect 212 429 227 446
rect 271 442 338 449
rect 7 419 80 420
rect 271 425 295 442
rect 312 425 338 442
rect 591 441 611 490
rect 646 463 655 490
rect 673 473 681 490
rect 672 463 681 473
rect 646 456 681 463
rect 21 385 123 402
rect 140 385 157 402
rect 174 385 191 402
rect 208 385 228 402
rect 271 399 338 425
rect 393 424 401 441
rect 418 424 435 441
rect 452 424 469 441
rect 486 424 611 441
rect 715 451 732 476
rect 715 409 732 434
rect 21 377 228 385
rect 272 395 337 399
rect 272 378 295 395
rect 312 378 337 395
rect 393 380 401 397
rect 418 380 435 397
rect 452 380 469 397
rect 486 380 501 397
rect 715 383 732 392
rect 21 127 58 377
rect 272 370 337 378
rect 415 344 474 380
rect 617 367 732 383
rect 617 350 715 367
rect 617 344 732 350
rect 115 325 732 344
rect 115 312 715 325
rect 115 283 132 312
rect 115 253 132 266
rect 159 283 176 295
rect 159 228 176 266
rect 215 283 232 312
rect 215 253 232 266
rect 259 283 276 295
rect 259 228 276 266
rect 315 283 332 312
rect 315 253 332 266
rect 359 283 376 295
rect 359 228 376 266
rect 415 283 432 312
rect 415 253 432 266
rect 459 283 476 295
rect 459 228 476 266
rect 515 283 532 312
rect 515 253 532 266
rect 559 283 576 295
rect 559 228 576 266
rect 615 283 632 312
rect 615 253 632 266
rect 659 283 676 295
rect 659 228 676 266
rect 715 283 732 308
rect 715 253 732 266
rect 759 451 776 476
rect 759 409 776 434
rect 759 367 776 392
rect 759 325 776 350
rect 759 283 776 308
rect 759 234 776 266
rect 817 355 834 527
rect 817 319 834 337
rect 817 283 834 301
rect 817 253 834 266
rect 861 348 878 361
rect 861 313 878 331
rect 861 277 878 295
rect 759 228 843 234
rect 99 211 117 228
rect 134 211 142 228
rect 159 211 217 228
rect 234 211 242 228
rect 259 211 317 228
rect 334 211 342 228
rect 359 211 417 228
rect 434 211 442 228
rect 459 211 517 228
rect 534 211 542 228
rect 559 211 617 228
rect 634 211 642 228
rect 659 211 717 228
rect 734 211 742 228
rect 759 211 792 228
rect 809 211 818 228
rect 835 211 843 228
rect 115 173 132 186
rect 115 127 132 156
rect 159 173 176 211
rect 159 144 176 156
rect 215 173 232 186
rect 215 127 232 156
rect 259 173 276 211
rect 259 144 276 156
rect 315 173 332 186
rect 315 127 332 156
rect 359 173 376 211
rect 359 144 376 156
rect 415 173 432 186
rect 415 127 432 156
rect 459 173 476 211
rect 459 144 476 156
rect 515 173 532 186
rect 515 127 532 156
rect 559 173 576 211
rect 559 144 576 156
rect 615 173 632 186
rect 615 127 632 156
rect 659 173 676 211
rect 759 205 843 211
rect 861 231 878 259
rect 861 208 902 231
rect 659 144 676 156
rect 715 173 732 186
rect 715 139 732 156
rect 700 127 715 133
rect 21 122 715 127
rect 21 105 732 122
rect 21 95 715 105
rect 700 90 715 95
rect 715 77 732 88
rect 759 173 776 205
rect 759 139 776 156
rect 817 167 834 187
rect 817 133 834 150
rect 861 167 878 208
rect 861 133 878 150
rect 759 105 776 122
rect 759 77 776 88
rect 0 15 12 32
rect 29 15 46 32
rect 63 15 80 32
rect 97 15 114 32
rect 131 15 148 32
rect 165 15 182 32
rect 199 15 216 32
rect 233 15 250 32
rect 267 15 284 32
rect 301 15 318 32
rect 335 15 352 32
rect 369 15 386 32
rect 403 15 420 32
rect 437 15 454 32
rect 471 15 488 32
rect 505 15 522 32
rect 539 15 556 32
rect 573 15 590 32
rect 607 15 624 32
rect 641 15 658 32
rect 675 15 692 32
rect 709 15 726 32
rect 743 15 760 32
rect 777 15 794 32
rect 811 15 828 32
rect 845 15 862 32
rect 879 15 902 32
<< viali >>
rect 12 605 29 622
rect 46 605 63 622
rect 80 605 97 622
rect 114 605 131 622
rect 148 605 165 622
rect 182 605 199 622
rect 216 605 233 622
rect 250 605 267 622
rect 284 605 301 622
rect 318 605 335 622
rect 352 605 369 622
rect 386 605 403 622
rect 420 605 437 622
rect 454 605 471 622
rect 488 605 505 622
rect 522 605 539 622
rect 556 605 573 622
rect 590 605 607 622
rect 624 605 636 622
rect 636 605 641 622
rect 658 605 675 622
rect 692 605 708 622
rect 708 605 709 622
rect 726 605 732 622
rect 732 605 743 622
rect 760 605 777 622
rect 794 605 804 622
rect 804 605 811 622
rect 828 605 845 622
rect 862 605 879 622
rect 25 506 42 523
rect 436 510 458 530
rect 591 524 608 529
rect 591 512 608 524
rect 711 539 728 556
rect 295 425 312 442
rect 655 473 672 480
rect 655 463 672 473
rect 295 378 312 395
rect 82 211 99 228
rect 792 211 809 228
rect 817 150 834 167
rect 12 15 29 32
rect 46 15 63 32
rect 80 15 97 32
rect 114 15 131 32
rect 148 15 165 32
rect 182 15 199 32
rect 216 15 233 32
rect 250 15 267 32
rect 284 15 301 32
rect 318 15 335 32
rect 352 15 369 32
rect 386 15 403 32
rect 420 15 437 32
rect 454 15 471 32
rect 488 15 505 32
rect 522 15 539 32
rect 556 15 573 32
rect 590 15 607 32
rect 624 15 641 32
rect 658 15 675 32
rect 692 15 709 32
rect 726 15 743 32
rect 760 15 777 32
rect 794 15 811 32
rect 828 15 845 32
rect 862 15 879 32
<< metal1 >>
rect 0 622 902 640
rect 0 605 12 622
rect 29 605 46 622
rect 63 605 80 622
rect 97 605 114 622
rect 131 605 148 622
rect 165 605 182 622
rect 199 605 216 622
rect 233 605 250 622
rect 267 605 284 622
rect 301 605 318 622
rect 335 605 352 622
rect 369 605 386 622
rect 403 605 420 622
rect 437 605 454 622
rect 471 605 488 622
rect 505 605 522 622
rect 539 605 556 622
rect 573 605 590 622
rect 607 605 624 622
rect 641 605 658 622
rect 675 605 692 622
rect 709 605 726 622
rect 743 605 760 622
rect 777 605 794 622
rect 811 605 828 622
rect 845 605 862 622
rect 879 605 902 622
rect 0 592 902 605
rect 705 556 734 562
rect 705 539 711 556
rect 728 539 734 556
rect 19 530 464 536
rect 705 534 734 539
rect 19 523 436 530
rect 19 506 25 523
rect 42 510 436 523
rect 458 510 464 530
rect 42 506 464 510
rect 585 529 735 534
rect 585 512 591 529
rect 608 512 735 529
rect 585 507 735 512
rect 19 500 464 506
rect 649 480 890 488
rect 649 463 655 480
rect 672 463 890 480
rect 649 457 890 463
rect 272 449 337 450
rect 271 442 338 449
rect 271 425 295 442
rect 312 425 338 442
rect 271 395 338 425
rect 271 378 295 395
rect 312 378 338 395
rect 271 345 338 378
rect 5 297 902 345
rect 76 228 813 234
rect 76 211 82 228
rect 99 211 792 228
rect 809 211 813 228
rect 76 206 813 211
rect 76 205 812 206
rect 871 173 891 297
rect 811 167 891 173
rect 811 150 817 167
rect 834 150 891 167
rect 811 144 891 150
rect 0 32 902 48
rect 0 15 12 32
rect 29 15 46 32
rect 63 15 80 32
rect 97 15 114 32
rect 131 15 148 32
rect 165 15 182 32
rect 199 15 216 32
rect 233 15 250 32
rect 267 15 284 32
rect 301 15 318 32
rect 335 15 352 32
rect 369 15 386 32
rect 403 15 420 32
rect 437 15 454 32
rect 471 15 488 32
rect 505 15 522 32
rect 539 15 556 32
rect 573 15 590 32
rect 607 15 624 32
rect 641 15 658 32
rect 675 15 692 32
rect 709 15 726 32
rect 743 15 760 32
rect 777 15 794 32
rect 811 15 828 32
rect 845 15 862 32
rect 879 15 902 32
rect 0 0 902 15
<< labels >>
rlabel locali 902 208 902 231 7 Clk_Out
port 5 w signal output
rlabel metal1 0 0 0 48 3 VDD
port 3 e power bidirectional
rlabel metal1 5 297 5 345 3 GND
port 4 e ground bidirectional
rlabel metal1 0 592 0 640 3 VDD
port 3 e power bidirectional
rlabel locali 7 419 7 439 3 VCtrl
port 2 e signal input
rlabel metal1 890 457 890 488 1 ENb
port 6 n signal input
<< properties >>
string LEFsite unithddb1
string LEFclass CORE
<< end >>
