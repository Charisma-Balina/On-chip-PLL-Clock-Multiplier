* SKY130 Spice File.
.param
+ tol_nfom = 0.069u
+ tol_pfom = 0.060u
+ tol_nw = 0.069u
+ tol_poly = 0.041u
+ tol_li = 0.020u
+ tol_m1 = 0.025u
+ tol_m2 = 0.025u
+ tol_m3 = 0.065u
+ tol_m4 = 0.065u
+ tol_m5 = 0.17u
+ tol_rdl = 1.0u
.param
+ rcn=70
+ rcp=330
+ rdn=108
+ rdp=166
+ rdn_hv=102
+ rdp_hv=160
+ rp1=42.2
+ rnw=1240
+ rl1=9.5
+ rm1= 0.105
+ rm2= 0.105
+ rm3= 0.038
+ rm4= 0.038
+ rm5= 0.0212
+ rrdl= 0.004
+ rcp1=25.28
+ rcl1=1.6
+ rcvia=2.0
+ rcvia2=0.50
+ rcvia3=0.50
+ rcvia4=0.012
+ rcrdlcon=0.0046
+ rspwres=2803
* P+ Poly Preres Parameters
.param
+ crpf_precision=  1.53e-04   $ Units: farad/meter^2
+ crpfsw_precision_1_1=  5.83e-11 $ Units: farad/meter
+ crpfsw_precision_2_1=  6.19e-11 $ Units: farad/meter
+ crpfsw_precision_4_1=  6.66e-11 $ Units: farad/meter
+ crpfsw_precision_8_2=  7.22e-11 $ Units: farad/meter
+ crpfsw_precision_16_2=  7.88e-11 $ Units: farad/meter
.include "../sky130_fd_pr__model__r+c.model.spice"
.include "../parameters/slow.spice"
