* SKY130 Spice File.
.param
+ tol_nfom = -0.0483u
+ tol_pfom = -0.042u
+ tol_nw = -0.0483u
+ tol_poly = -0.0287u
+ tol_li = -0.014u
+ tol_m1 = -0.0175u
+ tol_m2 = -0.0175u
+ tol_m3 = -0.0455u
+ tol_m4 = -0.0455u
+ tol_m5 = -0.119u
+ tol_rdl = -0.7u
.param
+ rcn=296.1
+ rcp=789
+ rdn=128.4
+ rdp=218.7
+ rdn_hv=122.4
+ rdp_hv=212.7
+ rp1=53.52
+ rnw=2022
+ rl1=14.02
+ rm1=0.139
+ rm2=0.139
+ rm3=0.0533
+ rm4=0.0533
+ rm5=0.03361
+ rrdl=0.00617
+ rcp1=213.88
+ rcl1=18.61
+ rcvia=11.85
+ rcvia2=6.623
+ rcvia3=6.623
+ rcvia4=0.7377
+ rcrdlcon=0.00713
+ rspwres=4120
* P+ Poly Preres Parameters
.param
+ crpf_precision=  1.39e-04   $ Units: farad/meter^2
+ crpfsw_precision_1_1=  5.59e-11 $ Units: farad/meter
+ crpfsw_precision_2_1=  5.95e-11 $ Units: farad/meter
+ crpfsw_precision_4_1=  6.41e-11 $ Units: farad/meter
+ crpfsw_precision_8_2=  6.96e-11 $ Units: farad/meter
+ crpfsw_precision_16_2=  7.61e-11 $ Units: farad/meter
.include "../sky130_fd_pr__model__r+c.model.spice"
.include "../parameters/slow_70p.spice"
