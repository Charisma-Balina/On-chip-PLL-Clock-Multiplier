* SKY130 Spice File.
* RF MOS Parameters
.include "../../../cells/rf_nfet_01v8/sky130_fd_pr__rf_nfet_01v8_b__sf.corner.spice"
.include "../../../cells/rf_nfet_01v8_lvt/sky130_fd_pr__rf_nfet_01v8_lvt_b__sf.corner.spice"
.include "../../../cells/rf_nfet_g5v0d10v5/sky130_fd_pr__rf_nfet_g5v0d10v5_b__sf.corner.spice"
.include "../../../cells/rf_pfet_01v8/sky130_fd_pr__rf_pfet_01v8_b__sf.corner.spice"
.include "../../../cells/rf_nfet_01v8/sky130_fd_pr__rf_nfet_01v8__mismatch.corner.spice"
.include "../../../cells/rf_nfet_01v8_lvt/sky130_fd_pr__rf_nfet_01v8_lvt__mismatch.corner.spice"
.include "../../../cells/rf_nfet_g5v0d10v5/sky130_fd_pr__rf_nfet_g5v0d10v5__mismatch.corner.spice"
.include "../../../cells/rf_pfet_01v8/sky130_fd_pr__rf_pfet_01v8__mismatch.corner.spice"
.include "../../../cells/rf_pfet_01v8_mvt/sky130_fd_pr__rf_pfet_01v8_mvt__sf_discrete.corner.spice"
.include "../../../cells/rf_pfet_01v8_mvt/sky130_fd_pr__rf_pfet_01v8_mvt__mismatch.corner.spice"
