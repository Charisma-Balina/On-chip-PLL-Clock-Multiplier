* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0

.SUBCKT sky130_fd_pr__pfet_01v8_aM04W1p65L0p18 BULK DRAIN GATE SOURCE
*.PININFO BULK:? DRAIN:? GATE:? SOURCE:?
M1 DRAIN GATE BULK model_use_only w=1.65 l=0.18 m=1
M2 DRAIN GATE BULK model_use_only w=1.65 l=0.18 m=1
M3 DRAIN GATE BULK model_use_only w=1.65 l=0.18 m=1
M4 DRAIN GATE BULK model_use_only w=1.65 l=0.18 m=1
.ENDS sky130_fd_pr__pfet_01v8_aM04W1p65L0p18
