* SKY130 Spice File.
* Slow    Varactor Parameters
.param
+ cnwvc_tox='41.6503*1.024*1.06'
+ cnwvc_cdepmult=0.9
+ cnwvc_cintmult=0.95
+ cnwvc_vt1='0.3333+0.112'
+ cnwvc_vt2='0.2380952+0.112'
+ cnwvc_vtr='0.16+0.112'
+ cnwvc_dwc=-0.02
+ cnwvc_dlc=-0.01
+ cnwvc_dld=-0.0008
+ cnwvc2_tox='41.7642*1.017*1.06'
+ cnwvc2_cdepmult=0.95
+ cnwvc2_cintmult=0.95
+ cnwvc2_vt1='0.2+0.074'
+ cnwvc2_vt2='0.33+0.074'
+ cnwvc2_vtr='0.14+0.074'
+ cnwvc2_dwc=-0.02
+ cnwvc2_dlc=-0.01
+ cnwvc2_dld=-0.0006
* sky130_fd_pr__model__parasitic__diode_ps2nw Parameters
.param
+ sky130_fd_pr__model__parasitic__diode_ps2nw__ajunction_mult = 7.9012e-01    $ Units: farad/meter^2
+ sky130_fd_pr__model__parasitic__diode_ps2nw__pjunction_mult = 9.1728e-01    $ Units: farad/meter^2
* sky130_fd_pr__model__parasitic__diode_ps2dn Parameters
+ sky130_fd_pr__model__parasitic__diode_ps2dn__ajunction_mult = 0.710       $ Units: farad/meter
+ sky130_fd_pr__model__parasitic__diode_ps2dn__pjunction_mult = 7.0406e-01  $ Units: farad/meter
* sky130_fd_pr__model__parasitic__diode_pw2dn Parameters
+ sky130_fd_pr__model__parasitic__diode_pw2dn__ajunction_mult = 0.69      $ Units: farad/meter
+ sky130_fd_pr__model__parasitic__diode_pw2dn__pjunction_mult = 8.7913e-01 $ Units: farad/meter
* sky130_fd_pr__diode_pw2nd_05v5  Parameters
+ sky130_fd_pr__nfet_01v8__ajunction_mult = 0.7739
+ sky130_fd_pr__nfet_01v8__pjunction_mult = 0.79336
* sky130_fd_pr__diode_pd2nw_05v5_hvt  Parameters
+ sky130_fd_pr__pfet_01v8_hvt__ajunction_mult = 1.0771e+0
+ sky130_fd_pr__pfet_01v8_hvt__pjunction_mult = 1.1263e+0
+ dkispp=9.2840e-01 dkbfpp=9.5154e-01 dknfpp=1.000
+ dkispp5x=1.0046e+00 dkbfpp5x=1.1288e+00 dknfpp5x=1.0009e+00 dkisepp5x=0.745
+ cvpp2_nhvnative10x4_cor=1.136
+ cvpp2_nhvnative10x4_sub=1.23e-14
+ cvpp2_phv5x4_cor=0.862
+ cvpp2_phv5x4_sub=8.68e-16
