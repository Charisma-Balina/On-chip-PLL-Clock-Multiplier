magic
tech sky130A
timestamp 1606013393
<< nwell >>
rect 12 252 171 297
rect 12 144 346 252
<< nmos >>
rect 65 74 80 110
rect 171 74 186 110
rect 284 74 299 110
<< pmos >>
rect 65 162 80 234
rect 171 162 186 234
rect 284 162 299 234
<< ndiff >>
rect 36 100 65 110
rect 36 83 42 100
rect 59 83 65 100
rect 36 74 65 83
rect 80 100 109 110
rect 80 83 86 100
rect 103 83 109 100
rect 80 74 109 83
rect 142 100 171 110
rect 142 83 148 100
rect 165 83 171 100
rect 142 74 171 83
rect 186 100 215 110
rect 186 83 192 100
rect 209 83 215 100
rect 186 74 215 83
rect 255 100 284 110
rect 255 83 261 100
rect 278 83 284 100
rect 255 74 284 83
rect 299 100 328 110
rect 299 83 305 100
rect 322 83 328 100
rect 299 74 328 83
<< pdiff >>
rect 36 225 65 234
rect 36 208 42 225
rect 59 208 65 225
rect 36 191 65 208
rect 36 174 42 191
rect 59 174 65 191
rect 36 162 65 174
rect 80 217 109 234
rect 80 200 86 217
rect 103 200 109 217
rect 80 183 109 200
rect 80 166 86 183
rect 103 166 109 183
rect 80 162 109 166
rect 142 217 171 234
rect 142 200 148 217
rect 165 200 171 217
rect 142 183 171 200
rect 142 166 148 183
rect 165 166 171 183
rect 142 162 171 166
rect 186 217 215 234
rect 186 200 192 217
rect 209 200 215 217
rect 186 183 215 200
rect 186 166 192 183
rect 209 166 215 183
rect 186 162 215 166
rect 255 217 284 234
rect 255 200 261 217
rect 278 200 284 217
rect 255 183 284 200
rect 255 166 261 183
rect 278 166 284 183
rect 255 162 284 166
rect 299 217 328 234
rect 299 200 305 217
rect 322 200 328 217
rect 299 183 328 200
rect 299 166 305 183
rect 322 166 328 183
rect 299 162 328 166
<< ndiffc >>
rect 42 83 59 100
rect 86 83 103 100
rect 148 83 165 100
rect 192 83 209 100
rect 261 83 278 100
rect 305 83 322 100
<< pdiffc >>
rect 42 208 59 225
rect 42 174 59 191
rect 86 200 103 217
rect 86 166 103 183
rect 148 200 165 217
rect 148 166 165 183
rect 192 200 209 217
rect 192 166 209 183
rect 261 200 278 217
rect 261 166 278 183
rect 305 200 322 217
rect 305 166 322 183
<< psubdiff >>
rect 30 1 42 18
rect 59 1 71 18
<< nsubdiff >>
rect 30 262 42 279
rect 59 262 71 279
<< psubdiffcont >>
rect 42 1 59 18
<< nsubdiffcont >>
rect 42 262 59 279
<< poly >>
rect 163 280 196 285
rect 163 263 171 280
rect 188 263 196 280
rect 163 258 196 263
rect 276 280 309 285
rect 276 263 284 280
rect 301 263 309 280
rect 276 258 309 263
rect 65 234 80 247
rect 171 234 186 258
rect 284 234 299 258
rect 65 110 80 162
rect 171 149 186 162
rect 284 149 299 162
rect 171 110 186 123
rect 284 110 299 123
rect 65 59 80 74
rect 171 59 186 74
rect 284 59 299 74
rect 65 54 110 59
rect 65 37 84 54
rect 101 37 110 54
rect 65 32 110 37
rect 163 54 196 59
rect 163 37 171 54
rect 188 37 196 54
rect 163 32 196 37
rect 276 54 309 59
rect 276 37 284 54
rect 301 37 309 54
rect 276 32 309 37
<< polycont >>
rect 171 263 188 280
rect 284 263 301 280
rect 84 37 101 54
rect 171 37 188 54
rect 284 37 301 54
<< locali >>
rect 42 279 59 293
rect 42 225 59 262
rect 42 191 59 208
rect 42 162 59 174
rect 86 280 244 282
rect 86 263 171 280
rect 188 263 244 280
rect 276 263 284 280
rect 301 263 309 280
rect 86 261 244 263
rect 86 217 103 261
rect 86 183 103 200
rect 42 100 59 110
rect 42 20 59 83
rect 86 100 103 166
rect 148 217 165 234
rect 148 183 165 200
rect 148 149 165 166
rect 133 143 165 149
rect 133 126 135 143
rect 152 126 165 143
rect 133 122 165 126
rect 86 74 103 83
rect 148 100 165 122
rect 148 74 165 83
rect 192 217 209 234
rect 192 183 209 200
rect 192 145 209 166
rect 192 100 209 128
rect 192 74 209 83
rect 227 57 244 261
rect 261 229 278 234
rect 261 183 278 200
rect 261 100 278 166
rect 261 74 278 83
rect 305 232 322 234
rect 305 229 334 232
rect 305 217 314 229
rect 331 212 334 229
rect 322 209 334 212
rect 305 183 322 200
rect 305 100 322 166
rect 305 74 322 83
rect 163 54 196 56
rect 76 37 84 54
rect 101 37 109 54
rect 163 37 171 54
rect 188 37 196 54
rect 163 35 196 37
rect 227 54 309 57
rect 227 37 284 54
rect 301 37 309 54
rect 227 36 309 37
rect 30 18 71 20
rect 30 1 42 18
rect 59 1 71 18
rect 30 0 71 1
<< viali >>
rect 284 263 301 280
rect 135 126 152 143
rect 192 128 209 145
rect 261 217 278 229
rect 261 212 278 217
rect 314 217 331 229
rect 314 212 322 217
rect 322 212 331 217
rect 84 37 101 54
rect 171 37 188 54
<< metal1 >>
rect 276 284 308 287
rect 276 258 279 284
rect 305 258 308 284
rect 276 255 308 258
rect 0 229 284 235
rect 0 212 261 229
rect 278 212 284 229
rect 0 206 284 212
rect 308 229 390 235
rect 308 212 314 229
rect 331 212 390 229
rect 308 206 390 212
rect 363 188 390 206
rect 363 151 408 188
rect 0 143 158 150
rect 0 126 135 143
rect 152 126 158 143
rect 0 120 158 126
rect 186 146 408 151
rect 186 145 392 146
rect 186 128 192 145
rect 209 128 392 145
rect 186 122 392 128
rect 163 60 195 61
rect 0 58 195 60
rect 0 54 166 58
rect 0 37 84 54
rect 101 37 166 54
rect 0 32 166 37
rect 192 32 195 58
rect 0 30 195 32
rect 163 29 195 30
<< via1 >>
rect 279 280 305 284
rect 279 263 284 280
rect 284 263 301 280
rect 301 263 305 280
rect 279 258 305 263
rect 166 54 192 58
rect 166 37 171 54
rect 171 37 188 54
rect 188 37 192 54
rect 166 32 192 37
<< metal2 >>
rect 276 284 308 287
rect 276 283 279 284
rect 223 258 279 283
rect 305 258 308 284
rect 163 60 195 61
rect 223 60 248 258
rect 276 255 308 258
rect 163 58 248 60
rect 163 32 166 58
rect 192 32 248 58
rect 163 30 248 32
rect 163 29 195 30
<< labels >>
rlabel metal1 0 30 0 60 3 SEL
port 1 e signal input
rlabel metal1 0 206 0 235 3 A
port 2 e signal input
rlabel metal1 0 120 0 150 3 B
port 3 e signal input
rlabel metal1 408 146 408 188 7 Out
port 4 w signal output
rlabel locali 42 12 59 12 1 GND
port 6 n power bidirectional
rlabel locali 42 293 59 293 5 VDD
port 5 s power bidirectional
<< properties >>
string LEFsite unithddb1
string LEFclass CORE
<< end >>
