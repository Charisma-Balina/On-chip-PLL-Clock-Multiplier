* SKY130 Spice File.
.param  globalk=1
.param  localkswitch=1
.param  capunits = '1.0*1e-6'
.param
+ mcp1f_ca_w_0_150_s_0_210 = 1.36e-04  mcp1f_cc_w_0_150_s_0_210 = 8.49e-11  mcp1f_cf_w_0_150_s_0_210 = 1.21e-11
+ mcp1f_ca_w_0_150_s_0_263 = 1.36e-04  mcp1f_cc_w_0_150_s_0_263 = 6.71e-11  mcp1f_cf_w_0_150_s_0_263 = 1.49e-11
+ mcp1f_ca_w_0_150_s_0_315 = 1.36e-04  mcp1f_cc_w_0_150_s_0_315 = 5.63e-11  mcp1f_cf_w_0_150_s_0_315 = 1.74e-11
+ mcp1f_ca_w_0_150_s_0_420 = 1.36e-04  mcp1f_cc_w_0_150_s_0_420 = 4.21e-11  mcp1f_cf_w_0_150_s_0_420 = 2.20e-11
+ mcp1f_ca_w_0_150_s_0_525 = 1.36e-04  mcp1f_cc_w_0_150_s_0_525 = 3.39e-11  mcp1f_cf_w_0_150_s_0_525 = 2.58e-11
+ mcp1f_ca_w_0_150_s_0_630 = 1.36e-04  mcp1f_cc_w_0_150_s_0_630 = 2.81e-11  mcp1f_cf_w_0_150_s_0_630 = 2.91e-11
+ mcp1f_ca_w_0_150_s_0_840 = 1.36e-04  mcp1f_cc_w_0_150_s_0_840 = 2.03e-11  mcp1f_cf_w_0_150_s_0_840 = 3.44e-11
+ mcp1f_ca_w_0_150_s_1_260 = 1.36e-04  mcp1f_cc_w_0_150_s_1_260 = 1.16e-11  mcp1f_cf_w_0_150_s_1_260 = 4.15e-11
+ mcp1f_ca_w_0_150_s_2_310 = 1.36e-04  mcp1f_cc_w_0_150_s_2_310 = 4.90e-12  mcp1f_cf_w_0_150_s_2_310 = 4.77e-11
+ mcp1f_ca_w_0_150_s_5_250 = 1.36e-04  mcp1f_cc_w_0_150_s_5_250 = 1.10e-12  mcp1f_cf_w_0_150_s_5_250 = 5.15e-11
+ mcp1f_ca_w_1_200_s_0_210 = 1.36e-04  mcp1f_cc_w_1_200_s_0_210 = 1.03e-10  mcp1f_cf_w_1_200_s_0_210 = 1.21e-11
+ mcp1f_ca_w_1_200_s_0_263 = 1.36e-04  mcp1f_cc_w_1_200_s_0_263 = 8.44e-11  mcp1f_cf_w_1_200_s_0_263 = 1.49e-11
+ mcp1f_ca_w_1_200_s_0_315 = 1.36e-04  mcp1f_cc_w_1_200_s_0_315 = 7.23e-11  mcp1f_cf_w_1_200_s_0_315 = 1.74e-11
+ mcp1f_ca_w_1_200_s_0_420 = 1.36e-04  mcp1f_cc_w_1_200_s_0_420 = 5.69e-11  mcp1f_cf_w_1_200_s_0_420 = 2.19e-11
+ mcp1f_ca_w_1_200_s_0_525 = 1.36e-04  mcp1f_cc_w_1_200_s_0_525 = 4.72e-11  mcp1f_cf_w_1_200_s_0_525 = 2.59e-11
+ mcp1f_ca_w_1_200_s_0_630 = 1.36e-04  mcp1f_cc_w_1_200_s_0_630 = 4.04e-11  mcp1f_cf_w_1_200_s_0_630 = 2.93e-11
+ mcp1f_ca_w_1_200_s_0_840 = 1.36e-04  mcp1f_cc_w_1_200_s_0_840 = 3.13e-11  mcp1f_cf_w_1_200_s_0_840 = 3.49e-11
+ mcp1f_ca_w_1_200_s_1_260 = 1.36e-04  mcp1f_cc_w_1_200_s_1_260 = 2.11e-11  mcp1f_cf_w_1_200_s_1_260 = 4.25e-11
+ mcp1f_ca_w_1_200_s_2_310 = 1.36e-04  mcp1f_cc_w_1_200_s_2_310 = 1.05e-11  mcp1f_cf_w_1_200_s_2_310 = 5.20e-11
+ mcp1f_ca_w_1_200_s_5_250 = 1.36e-04  mcp1f_cc_w_1_200_s_5_250 = 3.30e-12  mcp1f_cf_w_1_200_s_5_250 = 5.90e-11
+ mcl1f_ca_w_0_170_s_0_180 = 4.51e-05  mcl1f_cc_w_0_170_s_0_180 = 9.37e-11  mcl1f_cf_w_0_170_s_0_180 = 3.46e-12
+ mcl1f_ca_w_0_170_s_0_225 = 4.51e-05  mcl1f_cc_w_0_170_s_0_225 = 7.74e-11  mcl1f_cf_w_0_170_s_0_225 = 4.43e-12
+ mcl1f_ca_w_0_170_s_0_270 = 4.51e-05  mcl1f_cc_w_0_170_s_0_270 = 6.72e-11  mcl1f_cf_w_0_170_s_0_270 = 5.37e-12
+ mcl1f_ca_w_0_170_s_0_360 = 4.51e-05  mcl1f_cc_w_0_170_s_0_360 = 5.35e-11  mcl1f_cf_w_0_170_s_0_360 = 7.29e-12
+ mcl1f_ca_w_0_170_s_0_450 = 4.51e-05  mcl1f_cc_w_0_170_s_0_450 = 4.54e-11  mcl1f_cf_w_0_170_s_0_450 = 8.96e-12
+ mcl1f_ca_w_0_170_s_0_540 = 4.51e-05  mcl1f_cc_w_0_170_s_0_540 = 3.90e-11  mcl1f_cf_w_0_170_s_0_540 = 1.09e-11
+ mcl1f_ca_w_0_170_s_0_720 = 4.51e-05  mcl1f_cc_w_0_170_s_0_720 = 3.07e-11  mcl1f_cf_w_0_170_s_0_720 = 1.40e-11
+ mcl1f_ca_w_0_170_s_1_080 = 4.51e-05  mcl1f_cc_w_0_170_s_1_080 = 2.10e-11  mcl1f_cf_w_0_170_s_1_080 = 1.93e-11
+ mcl1f_ca_w_0_170_s_1_980 = 4.51e-05  mcl1f_cc_w_0_170_s_1_980 = 1.07e-11  mcl1f_cf_w_0_170_s_1_980 = 2.70e-11
+ mcl1f_ca_w_0_170_s_4_500 = 4.51e-05  mcl1f_cc_w_0_170_s_4_500 = 3.05e-12  mcl1f_cf_w_0_170_s_4_500 = 3.41e-11
+ mcl1f_ca_w_1_360_s_0_180 = 4.51e-05  mcl1f_cc_w_1_360_s_0_180 = 1.14e-10  mcl1f_cf_w_1_360_s_0_180 = 3.46e-12
+ mcl1f_ca_w_1_360_s_0_225 = 4.51e-05  mcl1f_cc_w_1_360_s_0_225 = 9.66e-11  mcl1f_cf_w_1_360_s_0_225 = 4.43e-12
+ mcl1f_ca_w_1_360_s_0_270 = 4.51e-05  mcl1f_cc_w_1_360_s_0_270 = 8.48e-11  mcl1f_cf_w_1_360_s_0_270 = 5.37e-12
+ mcl1f_ca_w_1_360_s_0_360 = 4.51e-05  mcl1f_cc_w_1_360_s_0_360 = 6.96e-11  mcl1f_cf_w_1_360_s_0_360 = 7.22e-12
+ mcl1f_ca_w_1_360_s_0_450 = 4.51e-05  mcl1f_cc_w_1_360_s_0_450 = 5.99e-11  mcl1f_cf_w_1_360_s_0_450 = 9.01e-12
+ mcl1f_ca_w_1_360_s_0_540 = 4.51e-05  mcl1f_cc_w_1_360_s_0_540 = 5.28e-11  mcl1f_cf_w_1_360_s_0_540 = 1.07e-11
+ mcl1f_ca_w_1_360_s_0_720 = 4.51e-05  mcl1f_cc_w_1_360_s_0_720 = 4.30e-11  mcl1f_cf_w_1_360_s_0_720 = 1.39e-11
+ mcl1f_ca_w_1_360_s_1_080 = 4.51e-05  mcl1f_cc_w_1_360_s_1_080 = 3.15e-11  mcl1f_cf_w_1_360_s_1_080 = 1.94e-11
+ mcl1f_ca_w_1_360_s_1_980 = 4.51e-05  mcl1f_cc_w_1_360_s_1_980 = 1.79e-11  mcl1f_cf_w_1_360_s_1_980 = 2.88e-11
+ mcl1f_ca_w_1_360_s_4_500 = 4.51e-05  mcl1f_cc_w_1_360_s_4_500 = 6.40e-12  mcl1f_cf_w_1_360_s_4_500 = 3.91e-11
+ mcl1d_ca_w_0_170_s_0_180 = 6.56e-05  mcl1d_cc_w_0_170_s_0_180 = 9.11e-11  mcl1d_cf_w_0_170_s_0_180 = 4.99e-12
+ mcl1d_ca_w_0_170_s_0_225 = 6.56e-05  mcl1d_cc_w_0_170_s_0_225 = 7.46e-11  mcl1d_cf_w_0_170_s_0_225 = 6.35e-12
+ mcl1d_ca_w_0_170_s_0_270 = 6.56e-05  mcl1d_cc_w_0_170_s_0_270 = 6.43e-11  mcl1d_cf_w_0_170_s_0_270 = 7.68e-12
+ mcl1d_ca_w_0_170_s_0_360 = 6.56e-05  mcl1d_cc_w_0_170_s_0_360 = 5.04e-11  mcl1d_cf_w_0_170_s_0_360 = 1.03e-11
+ mcl1d_ca_w_0_170_s_0_450 = 6.56e-05  mcl1d_cc_w_0_170_s_0_450 = 4.20e-11  mcl1d_cf_w_0_170_s_0_450 = 1.26e-11
+ mcl1d_ca_w_0_170_s_0_540 = 6.56e-05  mcl1d_cc_w_0_170_s_0_540 = 3.55e-11  mcl1d_cf_w_0_170_s_0_540 = 1.52e-11
+ mcl1d_ca_w_0_170_s_0_720 = 6.56e-05  mcl1d_cc_w_0_170_s_0_720 = 2.71e-11  mcl1d_cf_w_0_170_s_0_720 = 1.92e-11
+ mcl1d_ca_w_0_170_s_1_080 = 6.56e-05  mcl1d_cc_w_0_170_s_1_080 = 1.75e-11  mcl1d_cf_w_0_170_s_1_080 = 2.55e-11
+ mcl1d_ca_w_0_170_s_1_980 = 6.56e-05  mcl1d_cc_w_0_170_s_1_980 = 8.00e-12  mcl1d_cf_w_0_170_s_1_980 = 3.33e-11
+ mcl1d_ca_w_0_170_s_4_500 = 6.56e-05  mcl1d_cc_w_0_170_s_4_500 = 2.11e-12  mcl1d_cf_w_0_170_s_4_500 = 3.90e-11
+ mcl1d_ca_w_1_360_s_0_180 = 6.56e-05  mcl1d_cc_w_1_360_s_0_180 = 1.10e-10  mcl1d_cf_w_1_360_s_0_180 = 4.98e-12
+ mcl1d_ca_w_1_360_s_0_225 = 6.56e-05  mcl1d_cc_w_1_360_s_0_225 = 9.25e-11  mcl1d_cf_w_1_360_s_0_225 = 6.35e-12
+ mcl1d_ca_w_1_360_s_0_270 = 6.56e-05  mcl1d_cc_w_1_360_s_0_270 = 8.08e-11  mcl1d_cf_w_1_360_s_0_270 = 7.68e-12
+ mcl1d_ca_w_1_360_s_0_360 = 6.56e-05  mcl1d_cc_w_1_360_s_0_360 = 6.55e-11  mcl1d_cf_w_1_360_s_0_360 = 1.03e-11
+ mcl1d_ca_w_1_360_s_0_450 = 6.56e-05  mcl1d_cc_w_1_360_s_0_450 = 5.58e-11  mcl1d_cf_w_1_360_s_0_450 = 1.27e-11
+ mcl1d_ca_w_1_360_s_0_540 = 6.56e-05  mcl1d_cc_w_1_360_s_0_540 = 4.87e-11  mcl1d_cf_w_1_360_s_0_540 = 1.50e-11
+ mcl1d_ca_w_1_360_s_0_720 = 6.56e-05  mcl1d_cc_w_1_360_s_0_720 = 3.90e-11  mcl1d_cf_w_1_360_s_0_720 = 1.91e-11
+ mcl1d_ca_w_1_360_s_1_080 = 6.56e-05  mcl1d_cc_w_1_360_s_1_080 = 2.77e-11  mcl1d_cf_w_1_360_s_1_080 = 2.57e-11
+ mcl1d_ca_w_1_360_s_1_980 = 6.56e-05  mcl1d_cc_w_1_360_s_1_980 = 1.48e-11  mcl1d_cf_w_1_360_s_1_980 = 3.58e-11
+ mcl1d_ca_w_1_360_s_4_500 = 6.56e-05  mcl1d_cc_w_1_360_s_4_500 = 5.05e-12  mcl1d_cf_w_1_360_s_4_500 = 4.51e-11
+ mcl1p1_ca_w_0_170_s_0_180 = 1.40e-04  mcl1p1_cc_w_0_170_s_0_180 = 8.43e-11  mcl1p1_cf_w_0_170_s_0_180 = 1.03e-11
+ mcl1p1_ca_w_0_170_s_0_225 = 1.40e-04  mcl1p1_cc_w_0_170_s_0_225 = 6.78e-11  mcl1p1_cf_w_0_170_s_0_225 = 1.29e-11
+ mcl1p1_ca_w_0_170_s_0_270 = 1.40e-04  mcl1p1_cc_w_0_170_s_0_270 = 5.72e-11  mcl1p1_cf_w_0_170_s_0_270 = 1.55e-11
+ mcl1p1_ca_w_0_170_s_0_360 = 1.40e-04  mcl1p1_cc_w_0_170_s_0_360 = 4.30e-11  mcl1p1_cf_w_0_170_s_0_360 = 2.03e-11
+ mcl1p1_ca_w_0_170_s_0_450 = 1.40e-04  mcl1p1_cc_w_0_170_s_0_450 = 3.45e-11  mcl1p1_cf_w_0_170_s_0_450 = 2.41e-11
+ mcl1p1_ca_w_0_170_s_0_540 = 1.40e-04  mcl1p1_cc_w_0_170_s_0_540 = 2.78e-11  mcl1p1_cf_w_0_170_s_0_540 = 2.81e-11
+ mcl1p1_ca_w_0_170_s_0_720 = 1.40e-04  mcl1p1_cc_w_0_170_s_0_720 = 1.96e-11  mcl1p1_cf_w_0_170_s_0_720 = 3.37e-11
+ mcl1p1_ca_w_0_170_s_1_080 = 1.40e-04  mcl1p1_cc_w_0_170_s_1_080 = 1.12e-11  mcl1p1_cf_w_0_170_s_1_080 = 4.08e-11
+ mcl1p1_ca_w_0_170_s_1_980 = 1.40e-04  mcl1p1_cc_w_0_170_s_1_980 = 4.45e-12  mcl1p1_cf_w_0_170_s_1_980 = 4.71e-11
+ mcl1p1_ca_w_0_170_s_4_500 = 1.40e-04  mcl1p1_cc_w_0_170_s_4_500 = 1.10e-12  mcl1p1_cf_w_0_170_s_4_500 = 5.04e-11
+ mcl1p1_ca_w_1_360_s_0_180 = 1.40e-04  mcl1p1_cc_w_1_360_s_0_180 = 1.02e-10  mcl1p1_cf_w_1_360_s_0_180 = 1.04e-11
+ mcl1p1_ca_w_1_360_s_0_225 = 1.40e-04  mcl1p1_cc_w_1_360_s_0_225 = 8.45e-11  mcl1p1_cf_w_1_360_s_0_225 = 1.30e-11
+ mcl1p1_ca_w_1_360_s_0_270 = 1.40e-04  mcl1p1_cc_w_1_360_s_0_270 = 7.27e-11  mcl1p1_cf_w_1_360_s_0_270 = 1.55e-11
+ mcl1p1_ca_w_1_360_s_0_360 = 1.40e-04  mcl1p1_cc_w_1_360_s_0_360 = 5.75e-11  mcl1p1_cf_w_1_360_s_0_360 = 2.02e-11
+ mcl1p1_ca_w_1_360_s_0_450 = 1.40e-04  mcl1p1_cc_w_1_360_s_0_450 = 4.78e-11  mcl1p1_cf_w_1_360_s_0_450 = 2.43e-11
+ mcl1p1_ca_w_1_360_s_0_540 = 1.40e-04  mcl1p1_cc_w_1_360_s_0_540 = 4.09e-11  mcl1p1_cf_w_1_360_s_0_540 = 2.80e-11
+ mcl1p1_ca_w_1_360_s_0_720 = 1.40e-04  mcl1p1_cc_w_1_360_s_0_720 = 3.16e-11  mcl1p1_cf_w_1_360_s_0_720 = 3.39e-11
+ mcl1p1_ca_w_1_360_s_1_080 = 1.40e-04  mcl1p1_cc_w_1_360_s_1_080 = 2.12e-11  mcl1p1_cf_w_1_360_s_1_080 = 4.20e-11
+ mcl1p1_ca_w_1_360_s_1_980 = 1.40e-04  mcl1p1_cc_w_1_360_s_1_980 = 1.05e-11  mcl1p1_cf_w_1_360_s_1_980 = 5.17e-11
+ mcl1p1_ca_w_1_360_s_4_500 = 1.40e-04  mcl1p1_cc_w_1_360_s_4_500 = 3.45e-12  mcl1p1_cf_w_1_360_s_4_500 = 5.87e-11
+ mcm1f_ca_w_0_140_s_0_140 = 3.18e-05  mcm1f_cc_w_0_140_s_0_140 = 1.22e-10  mcm1f_cf_w_0_140_s_0_140 = 1.86e-12
+ mcm1f_ca_w_0_140_s_0_175 = 3.18e-05  mcm1f_cc_w_0_140_s_0_175 = 1.17e-10  mcm1f_cf_w_0_140_s_0_175 = 2.41e-12
+ mcm1f_ca_w_0_140_s_0_210 = 3.18e-05  mcm1f_cc_w_0_140_s_0_210 = 1.11e-10  mcm1f_cf_w_0_140_s_0_210 = 2.97e-12
+ mcm1f_ca_w_0_140_s_0_280 = 3.18e-05  mcm1f_cc_w_0_140_s_0_280 = 9.64e-11  mcm1f_cf_w_0_140_s_0_280 = 4.05e-12
+ mcm1f_ca_w_0_140_s_0_350 = 3.18e-05  mcm1f_cc_w_0_140_s_0_350 = 8.24e-11  mcm1f_cf_w_0_140_s_0_350 = 5.11e-12
+ mcm1f_ca_w_0_140_s_0_420 = 3.18e-05  mcm1f_cc_w_0_140_s_0_420 = 7.19e-11  mcm1f_cf_w_0_140_s_0_420 = 6.18e-12
+ mcm1f_ca_w_0_140_s_0_560 = 3.18e-05  mcm1f_cc_w_0_140_s_0_560 = 5.73e-11  mcm1f_cf_w_0_140_s_0_560 = 8.13e-12
+ mcm1f_ca_w_0_140_s_0_840 = 3.18e-05  mcm1f_cc_w_0_140_s_0_840 = 4.14e-11  mcm1f_cf_w_0_140_s_0_840 = 1.18e-11
+ mcm1f_ca_w_0_140_s_1_540 = 3.18e-05  mcm1f_cc_w_0_140_s_1_540 = 2.42e-11  mcm1f_cf_w_0_140_s_1_540 = 1.95e-11
+ mcm1f_ca_w_0_140_s_3_500 = 3.18e-05  mcm1f_cc_w_0_140_s_3_500 = 9.21e-12  mcm1f_cf_w_0_140_s_3_500 = 3.08e-11
+ mcm1f_ca_w_1_120_s_0_140 = 3.18e-05  mcm1f_cc_w_1_120_s_0_140 = 1.47e-10  mcm1f_cf_w_1_120_s_0_140 = 1.92e-12
+ mcm1f_ca_w_1_120_s_0_175 = 3.18e-05  mcm1f_cc_w_1_120_s_0_175 = 1.40e-10  mcm1f_cf_w_1_120_s_0_175 = 2.47e-12
+ mcm1f_ca_w_1_120_s_0_210 = 3.18e-05  mcm1f_cc_w_1_120_s_0_210 = 1.33e-10  mcm1f_cf_w_1_120_s_0_210 = 3.02e-12
+ mcm1f_ca_w_1_120_s_0_280 = 3.18e-05  mcm1f_cc_w_1_120_s_0_280 = 1.15e-10  mcm1f_cf_w_1_120_s_0_280 = 4.10e-12
+ mcm1f_ca_w_1_120_s_0_350 = 3.18e-05  mcm1f_cc_w_1_120_s_0_350 = 1.00e-10  mcm1f_cf_w_1_120_s_0_350 = 5.16e-12
+ mcm1f_ca_w_1_120_s_0_420 = 3.18e-05  mcm1f_cc_w_1_120_s_0_420 = 8.79e-11  mcm1f_cf_w_1_120_s_0_420 = 6.21e-12
+ mcm1f_ca_w_1_120_s_0_560 = 3.18e-05  mcm1f_cc_w_1_120_s_0_560 = 7.08e-11  mcm1f_cf_w_1_120_s_0_560 = 8.23e-12
+ mcm1f_ca_w_1_120_s_0_840 = 3.18e-05  mcm1f_cc_w_1_120_s_0_840 = 5.22e-11  mcm1f_cf_w_1_120_s_0_840 = 1.20e-11
+ mcm1f_ca_w_1_120_s_1_540 = 3.18e-05  mcm1f_cc_w_1_120_s_1_540 = 3.20e-11  mcm1f_cf_w_1_120_s_1_540 = 1.99e-11
+ mcm1f_ca_w_1_120_s_3_500 = 3.18e-05  mcm1f_cc_w_1_120_s_3_500 = 1.37e-11  mcm1f_cf_w_1_120_s_3_500 = 3.27e-11
+ mcm1d_ca_w_0_140_s_0_140 = 4.07e-05  mcm1d_cc_w_0_140_s_0_140 = 1.21e-10  mcm1d_cf_w_0_140_s_0_140 = 2.38e-12
+ mcm1d_ca_w_0_140_s_0_175 = 4.07e-05  mcm1d_cc_w_0_140_s_0_175 = 1.15e-10  mcm1d_cf_w_0_140_s_0_175 = 3.09e-12
+ mcm1d_ca_w_0_140_s_0_210 = 4.07e-05  mcm1d_cc_w_0_140_s_0_210 = 1.09e-10  mcm1d_cf_w_0_140_s_0_210 = 3.79e-12
+ mcm1d_ca_w_0_140_s_0_280 = 4.07e-05  mcm1d_cc_w_0_140_s_0_280 = 9.51e-11  mcm1d_cf_w_0_140_s_0_280 = 5.17e-12
+ mcm1d_ca_w_0_140_s_0_350 = 4.07e-05  mcm1d_cc_w_0_140_s_0_350 = 8.09e-11  mcm1d_cf_w_0_140_s_0_350 = 6.51e-12
+ mcm1d_ca_w_0_140_s_0_420 = 4.07e-05  mcm1d_cc_w_0_140_s_0_420 = 7.01e-11  mcm1d_cf_w_0_140_s_0_420 = 7.86e-12
+ mcm1d_ca_w_0_140_s_0_560 = 4.07e-05  mcm1d_cc_w_0_140_s_0_560 = 5.54e-11  mcm1d_cf_w_0_140_s_0_560 = 1.03e-11
+ mcm1d_ca_w_0_140_s_0_840 = 4.07e-05  mcm1d_cc_w_0_140_s_0_840 = 3.92e-11  mcm1d_cf_w_0_140_s_0_840 = 1.48e-11
+ mcm1d_ca_w_0_140_s_1_540 = 4.07e-05  mcm1d_cc_w_0_140_s_1_540 = 2.19e-11  mcm1d_cf_w_0_140_s_1_540 = 2.37e-11
+ mcm1d_ca_w_0_140_s_3_500 = 4.07e-05  mcm1d_cc_w_0_140_s_3_500 = 7.66e-12  mcm1d_cf_w_0_140_s_3_500 = 3.52e-11
+ mcm1d_ca_w_1_120_s_0_140 = 4.07e-05  mcm1d_cc_w_1_120_s_0_140 = 1.44e-10  mcm1d_cf_w_1_120_s_0_140 = 2.46e-12
+ mcm1d_ca_w_1_120_s_0_175 = 4.07e-05  mcm1d_cc_w_1_120_s_0_175 = 1.37e-10  mcm1d_cf_w_1_120_s_0_175 = 3.17e-12
+ mcm1d_ca_w_1_120_s_0_210 = 4.07e-05  mcm1d_cc_w_1_120_s_0_210 = 1.29e-10  mcm1d_cf_w_1_120_s_0_210 = 3.88e-12
+ mcm1d_ca_w_1_120_s_0_280 = 4.07e-05  mcm1d_cc_w_1_120_s_0_280 = 1.12e-10  mcm1d_cf_w_1_120_s_0_280 = 5.25e-12
+ mcm1d_ca_w_1_120_s_0_350 = 4.07e-05  mcm1d_cc_w_1_120_s_0_350 = 9.76e-11  mcm1d_cf_w_1_120_s_0_350 = 6.60e-12
+ mcm1d_ca_w_1_120_s_0_420 = 4.07e-05  mcm1d_cc_w_1_120_s_0_420 = 8.52e-11  mcm1d_cf_w_1_120_s_0_420 = 7.92e-12
+ mcm1d_ca_w_1_120_s_0_560 = 4.07e-05  mcm1d_cc_w_1_120_s_0_560 = 6.80e-11  mcm1d_cf_w_1_120_s_0_560 = 1.04e-11
+ mcm1d_ca_w_1_120_s_0_840 = 4.07e-05  mcm1d_cc_w_1_120_s_0_840 = 4.95e-11  mcm1d_cf_w_1_120_s_0_840 = 1.50e-11
+ mcm1d_ca_w_1_120_s_1_540 = 4.07e-05  mcm1d_cc_w_1_120_s_1_540 = 2.94e-11  mcm1d_cf_w_1_120_s_1_540 = 2.41e-11
+ mcm1d_ca_w_1_120_s_3_500 = 4.07e-05  mcm1d_cc_w_1_120_s_3_500 = 1.19e-11  mcm1d_cf_w_1_120_s_3_500 = 3.74e-11
+ mcm1p1_ca_w_0_140_s_0_140 = 6.07e-05  mcm1p1_cc_w_0_140_s_0_140 = 1.19e-10  mcm1p1_cf_w_0_140_s_0_140 = 3.54e-12
+ mcm1p1_ca_w_0_140_s_0_175 = 6.07e-05  mcm1p1_cc_w_0_140_s_0_175 = 1.13e-10  mcm1p1_cf_w_0_140_s_0_175 = 4.59e-12
+ mcm1p1_ca_w_0_140_s_0_210 = 6.07e-05  mcm1p1_cc_w_0_140_s_0_210 = 1.07e-10  mcm1p1_cf_w_0_140_s_0_210 = 5.63e-12
+ mcm1p1_ca_w_0_140_s_0_280 = 6.07e-05  mcm1p1_cc_w_0_140_s_0_280 = 9.22e-11  mcm1p1_cf_w_0_140_s_0_280 = 7.66e-12
+ mcm1p1_ca_w_0_140_s_0_350 = 6.07e-05  mcm1p1_cc_w_0_140_s_0_350 = 7.77e-11  mcm1p1_cf_w_0_140_s_0_350 = 9.60e-12
+ mcm1p1_ca_w_0_140_s_0_420 = 6.07e-05  mcm1p1_cc_w_0_140_s_0_420 = 6.70e-11  mcm1p1_cf_w_0_140_s_0_420 = 1.15e-11
+ mcm1p1_ca_w_0_140_s_0_560 = 6.07e-05  mcm1p1_cc_w_0_140_s_0_560 = 5.16e-11  mcm1p1_cf_w_0_140_s_0_560 = 1.50e-11
+ mcm1p1_ca_w_0_140_s_0_840 = 6.07e-05  mcm1p1_cc_w_0_140_s_0_840 = 3.53e-11  mcm1p1_cf_w_0_140_s_0_840 = 2.10e-11
+ mcm1p1_ca_w_0_140_s_1_540 = 6.07e-05  mcm1p1_cc_w_0_140_s_1_540 = 1.82e-11  mcm1p1_cf_w_0_140_s_1_540 = 3.16e-11
+ mcm1p1_ca_w_0_140_s_3_500 = 6.07e-05  mcm1p1_cc_w_0_140_s_3_500 = 5.70e-12  mcm1p1_cf_w_0_140_s_3_500 = 4.26e-11
+ mcm1p1_ca_w_1_120_s_0_140 = 6.07e-05  mcm1p1_cc_w_1_120_s_0_140 = 1.40e-10  mcm1p1_cf_w_1_120_s_0_140 = 3.73e-12
+ mcm1p1_ca_w_1_120_s_0_175 = 6.07e-05  mcm1p1_cc_w_1_120_s_0_175 = 1.33e-10  mcm1p1_cf_w_1_120_s_0_175 = 4.77e-12
+ mcm1p1_ca_w_1_120_s_0_210 = 6.07e-05  mcm1p1_cc_w_1_120_s_0_210 = 1.25e-10  mcm1p1_cf_w_1_120_s_0_210 = 5.80e-12
+ mcm1p1_ca_w_1_120_s_0_280 = 6.07e-05  mcm1p1_cc_w_1_120_s_0_280 = 1.08e-10  mcm1p1_cf_w_1_120_s_0_280 = 7.82e-12
+ mcm1p1_ca_w_1_120_s_0_350 = 6.07e-05  mcm1p1_cc_w_1_120_s_0_350 = 9.29e-11  mcm1p1_cf_w_1_120_s_0_350 = 9.77e-12
+ mcm1p1_ca_w_1_120_s_0_420 = 6.07e-05  mcm1p1_cc_w_1_120_s_0_420 = 8.04e-11  mcm1p1_cf_w_1_120_s_0_420 = 1.16e-11
+ mcm1p1_ca_w_1_120_s_0_560 = 6.07e-05  mcm1p1_cc_w_1_120_s_0_560 = 6.34e-11  mcm1p1_cf_w_1_120_s_0_560 = 1.52e-11
+ mcm1p1_ca_w_1_120_s_0_840 = 6.07e-05  mcm1p1_cc_w_1_120_s_0_840 = 4.49e-11  mcm1p1_cf_w_1_120_s_0_840 = 2.13e-11
+ mcm1p1_ca_w_1_120_s_1_540 = 6.07e-05  mcm1p1_cc_w_1_120_s_1_540 = 2.55e-11  mcm1p1_cf_w_1_120_s_1_540 = 3.23e-11
+ mcm1p1_ca_w_1_120_s_3_500 = 6.07e-05  mcm1p1_cc_w_1_120_s_3_500 = 9.65e-12  mcm1p1_cf_w_1_120_s_3_500 = 4.56e-11
+ mcm1l1_ca_w_0_140_s_0_140 = 1.63e-04  mcm1l1_cc_w_0_140_s_0_140 = 1.09e-10  mcm1l1_cf_w_0_140_s_0_140 = 8.86e-12
+ mcm1l1_ca_w_0_140_s_0_175 = 1.63e-04  mcm1l1_cc_w_0_140_s_0_175 = 1.04e-10  mcm1l1_cf_w_0_140_s_0_175 = 1.17e-11
+ mcm1l1_ca_w_0_140_s_0_210 = 1.63e-04  mcm1l1_cc_w_0_140_s_0_210 = 9.83e-11  mcm1l1_cf_w_0_140_s_0_210 = 1.43e-11
+ mcm1l1_ca_w_0_140_s_0_280 = 1.63e-04  mcm1l1_cc_w_0_140_s_0_280 = 8.24e-11  mcm1l1_cf_w_0_140_s_0_280 = 1.93e-11
+ mcm1l1_ca_w_0_140_s_0_350 = 1.63e-04  mcm1l1_cc_w_0_140_s_0_350 = 6.80e-11  mcm1l1_cf_w_0_140_s_0_350 = 2.37e-11
+ mcm1l1_ca_w_0_140_s_0_420 = 1.63e-04  mcm1l1_cc_w_0_140_s_0_420 = 5.68e-11  mcm1l1_cf_w_0_140_s_0_420 = 2.78e-11
+ mcm1l1_ca_w_0_140_s_0_560 = 1.63e-04  mcm1l1_cc_w_0_140_s_0_560 = 4.19e-11  mcm1l1_cf_w_0_140_s_0_560 = 3.45e-11
+ mcm1l1_ca_w_0_140_s_0_840 = 1.63e-04  mcm1l1_cc_w_0_140_s_0_840 = 2.64e-11  mcm1l1_cf_w_0_140_s_0_840 = 4.41e-11
+ mcm1l1_ca_w_0_140_s_1_540 = 1.63e-04  mcm1l1_cc_w_0_140_s_1_540 = 1.18e-11  mcm1l1_cf_w_0_140_s_1_540 = 5.66e-11
+ mcm1l1_ca_w_0_140_s_3_500 = 1.63e-04  mcm1l1_cc_w_0_140_s_3_500 = 3.25e-12  mcm1l1_cf_w_0_140_s_3_500 = 6.53e-11
+ mcm1l1_ca_w_1_120_s_0_140 = 1.63e-04  mcm1l1_cc_w_1_120_s_0_140 = 1.28e-10  mcm1l1_cf_w_1_120_s_0_140 = 9.03e-12
+ mcm1l1_ca_w_1_120_s_0_175 = 1.63e-04  mcm1l1_cc_w_1_120_s_0_175 = 1.21e-10  mcm1l1_cf_w_1_120_s_0_175 = 1.18e-11
+ mcm1l1_ca_w_1_120_s_0_210 = 1.63e-04  mcm1l1_cc_w_1_120_s_0_210 = 1.13e-10  mcm1l1_cf_w_1_120_s_0_210 = 1.45e-11
+ mcm1l1_ca_w_1_120_s_0_280 = 1.63e-04  mcm1l1_cc_w_1_120_s_0_280 = 9.62e-11  mcm1l1_cf_w_1_120_s_0_280 = 1.94e-11
+ mcm1l1_ca_w_1_120_s_0_350 = 1.63e-04  mcm1l1_cc_w_1_120_s_0_350 = 8.11e-11  mcm1l1_cf_w_1_120_s_0_350 = 2.39e-11
+ mcm1l1_ca_w_1_120_s_0_420 = 1.63e-04  mcm1l1_cc_w_1_120_s_0_420 = 6.92e-11  mcm1l1_cf_w_1_120_s_0_420 = 2.79e-11
+ mcm1l1_ca_w_1_120_s_0_560 = 1.63e-04  mcm1l1_cc_w_1_120_s_0_560 = 5.29e-11  mcm1l1_cf_w_1_120_s_0_560 = 3.46e-11
+ mcm1l1_ca_w_1_120_s_0_840 = 1.63e-04  mcm1l1_cc_w_1_120_s_0_840 = 3.58e-11  mcm1l1_cf_w_1_120_s_0_840 = 4.45e-11
+ mcm1l1_ca_w_1_120_s_1_540 = 1.63e-04  mcm1l1_cc_w_1_120_s_1_540 = 1.88e-11  mcm1l1_cf_w_1_120_s_1_540 = 5.78e-11
+ mcm1l1_ca_w_1_120_s_3_500 = 1.63e-04  mcm1l1_cc_w_1_120_s_3_500 = 6.65e-12  mcm1l1_cf_w_1_120_s_3_500 = 6.96e-11
+ mcm2f_ca_w_0_140_s_0_140 = 2.13e-05  mcm2f_cc_w_0_140_s_0_140 = 1.23e-10  mcm2f_cf_w_0_140_s_0_140 = 1.26e-12
+ mcm2f_ca_w_0_140_s_0_175 = 2.13e-05  mcm2f_cc_w_0_140_s_0_175 = 1.18e-10  mcm2f_cf_w_0_140_s_0_175 = 1.62e-12
+ mcm2f_ca_w_0_140_s_0_210 = 2.13e-05  mcm2f_cc_w_0_140_s_0_210 = 1.12e-10  mcm2f_cf_w_0_140_s_0_210 = 1.99e-12
+ mcm2f_ca_w_0_140_s_0_280 = 2.13e-05  mcm2f_cc_w_0_140_s_0_280 = 9.70e-11  mcm2f_cf_w_0_140_s_0_280 = 2.73e-12
+ mcm2f_ca_w_0_140_s_0_350 = 2.13e-05  mcm2f_cc_w_0_140_s_0_350 = 8.39e-11  mcm2f_cf_w_0_140_s_0_350 = 3.44e-12
+ mcm2f_ca_w_0_140_s_0_420 = 2.13e-05  mcm2f_cc_w_0_140_s_0_420 = 7.36e-11  mcm2f_cf_w_0_140_s_0_420 = 4.19e-12
+ mcm2f_ca_w_0_140_s_0_560 = 2.13e-05  mcm2f_cc_w_0_140_s_0_560 = 5.91e-11  mcm2f_cf_w_0_140_s_0_560 = 5.53e-12
+ mcm2f_ca_w_0_140_s_0_840 = 2.13e-05  mcm2f_cc_w_0_140_s_0_840 = 4.37e-11  mcm2f_cf_w_0_140_s_0_840 = 8.16e-12
+ mcm2f_ca_w_0_140_s_1_540 = 2.13e-05  mcm2f_cc_w_0_140_s_1_540 = 2.72e-11  mcm2f_cf_w_0_140_s_1_540 = 1.39e-11
+ mcm2f_ca_w_0_140_s_3_500 = 2.13e-05  mcm2f_cc_w_0_140_s_3_500 = 1.19e-11  mcm2f_cf_w_0_140_s_3_500 = 2.40e-11
+ mcm2f_ca_w_1_120_s_0_140 = 2.13e-05  mcm2f_cc_w_1_120_s_0_140 = 1.50e-10  mcm2f_cf_w_1_120_s_0_140 = 1.29e-12
+ mcm2f_ca_w_1_120_s_0_175 = 2.13e-05  mcm2f_cc_w_1_120_s_0_175 = 1.43e-10  mcm2f_cf_w_1_120_s_0_175 = 1.65e-12
+ mcm2f_ca_w_1_120_s_0_210 = 2.13e-05  mcm2f_cc_w_1_120_s_0_210 = 1.35e-10  mcm2f_cf_w_1_120_s_0_210 = 2.02e-12
+ mcm2f_ca_w_1_120_s_0_280 = 2.13e-05  mcm2f_cc_w_1_120_s_0_280 = 1.18e-10  mcm2f_cf_w_1_120_s_0_280 = 2.75e-12
+ mcm2f_ca_w_1_120_s_0_350 = 2.13e-05  mcm2f_cc_w_1_120_s_0_350 = 1.03e-10  mcm2f_cf_w_1_120_s_0_350 = 3.48e-12
+ mcm2f_ca_w_1_120_s_0_420 = 2.13e-05  mcm2f_cc_w_1_120_s_0_420 = 9.09e-11  mcm2f_cf_w_1_120_s_0_420 = 4.20e-12
+ mcm2f_ca_w_1_120_s_0_560 = 2.13e-05  mcm2f_cc_w_1_120_s_0_560 = 7.36e-11  mcm2f_cf_w_1_120_s_0_560 = 5.58e-12
+ mcm2f_ca_w_1_120_s_0_840 = 2.13e-05  mcm2f_cc_w_1_120_s_0_840 = 5.54e-11  mcm2f_cf_w_1_120_s_0_840 = 8.25e-12
+ mcm2f_ca_w_1_120_s_1_540 = 2.13e-05  mcm2f_cc_w_1_120_s_1_540 = 3.55e-11  mcm2f_cf_w_1_120_s_1_540 = 1.41e-11
+ mcm2f_ca_w_1_120_s_3_500 = 2.13e-05  mcm2f_cc_w_1_120_s_3_500 = 1.68e-11  mcm2f_cf_w_1_120_s_3_500 = 2.53e-11
+ mcm2d_ca_w_0_140_s_0_140 = 2.49e-05  mcm2d_cc_w_0_140_s_0_140 = 1.23e-10  mcm2d_cf_w_0_140_s_0_140 = 1.47e-12
+ mcm2d_ca_w_0_140_s_0_175 = 2.49e-05  mcm2d_cc_w_0_140_s_0_175 = 1.17e-10  mcm2d_cf_w_0_140_s_0_175 = 1.90e-12
+ mcm2d_ca_w_0_140_s_0_210 = 2.49e-05  mcm2d_cc_w_0_140_s_0_210 = 1.11e-10  mcm2d_cf_w_0_140_s_0_210 = 2.34e-12
+ mcm2d_ca_w_0_140_s_0_280 = 2.49e-05  mcm2d_cc_w_0_140_s_0_280 = 9.60e-11  mcm2d_cf_w_0_140_s_0_280 = 3.19e-12
+ mcm2d_ca_w_0_140_s_0_350 = 2.49e-05  mcm2d_cc_w_0_140_s_0_350 = 8.33e-11  mcm2d_cf_w_0_140_s_0_350 = 4.03e-12
+ mcm2d_ca_w_0_140_s_0_420 = 2.49e-05  mcm2d_cc_w_0_140_s_0_420 = 7.29e-11  mcm2d_cf_w_0_140_s_0_420 = 4.89e-12
+ mcm2d_ca_w_0_140_s_0_560 = 2.49e-05  mcm2d_cc_w_0_140_s_0_560 = 5.82e-11  mcm2d_cf_w_0_140_s_0_560 = 6.46e-12
+ mcm2d_ca_w_0_140_s_0_840 = 2.49e-05  mcm2d_cc_w_0_140_s_0_840 = 4.26e-11  mcm2d_cf_w_0_140_s_0_840 = 9.48e-12
+ mcm2d_ca_w_0_140_s_1_540 = 2.49e-05  mcm2d_cc_w_0_140_s_1_540 = 2.58e-11  mcm2d_cf_w_0_140_s_1_540 = 1.59e-11
+ mcm2d_ca_w_0_140_s_3_500 = 2.49e-05  mcm2d_cc_w_0_140_s_3_500 = 1.07e-11  mcm2d_cf_w_0_140_s_3_500 = 2.65e-11
+ mcm2d_ca_w_1_120_s_0_140 = 2.49e-05  mcm2d_cc_w_1_120_s_0_140 = 1.48e-10  mcm2d_cf_w_1_120_s_0_140 = 1.51e-12
+ mcm2d_ca_w_1_120_s_0_175 = 2.49e-05  mcm2d_cc_w_1_120_s_0_175 = 1.41e-10  mcm2d_cf_w_1_120_s_0_175 = 1.94e-12
+ mcm2d_ca_w_1_120_s_0_210 = 2.49e-05  mcm2d_cc_w_1_120_s_0_210 = 1.34e-10  mcm2d_cf_w_1_120_s_0_210 = 2.37e-12
+ mcm2d_ca_w_1_120_s_0_280 = 2.49e-05  mcm2d_cc_w_1_120_s_0_280 = 1.16e-10  mcm2d_cf_w_1_120_s_0_280 = 3.23e-12
+ mcm2d_ca_w_1_120_s_0_350 = 2.49e-05  mcm2d_cc_w_1_120_s_0_350 = 1.01e-10  mcm2d_cf_w_1_120_s_0_350 = 4.07e-12
+ mcm2d_ca_w_1_120_s_0_420 = 2.49e-05  mcm2d_cc_w_1_120_s_0_420 = 8.91e-11  mcm2d_cf_w_1_120_s_0_420 = 4.90e-12
+ mcm2d_ca_w_1_120_s_0_560 = 2.49e-05  mcm2d_cc_w_1_120_s_0_560 = 7.21e-11  mcm2d_cf_w_1_120_s_0_560 = 6.51e-12
+ mcm2d_ca_w_1_120_s_0_840 = 2.49e-05  mcm2d_cc_w_1_120_s_0_840 = 5.37e-11  mcm2d_cf_w_1_120_s_0_840 = 9.59e-12
+ mcm2d_ca_w_1_120_s_1_540 = 2.49e-05  mcm2d_cc_w_1_120_s_1_540 = 3.38e-11  mcm2d_cf_w_1_120_s_1_540 = 1.62e-11
+ mcm2d_ca_w_1_120_s_3_500 = 2.49e-05  mcm2d_cc_w_1_120_s_3_500 = 1.54e-11  mcm2d_cf_w_1_120_s_3_500 = 2.81e-11
+ mcm2p1_ca_w_0_140_s_0_140 = 3.12e-05  mcm2p1_cc_w_0_140_s_0_140 = 1.22e-10  mcm2p1_cf_w_0_140_s_0_140 = 1.84e-12
+ mcm2p1_ca_w_0_140_s_0_175 = 3.12e-05  mcm2p1_cc_w_0_140_s_0_175 = 1.17e-10  mcm2p1_cf_w_0_140_s_0_175 = 2.38e-12
+ mcm2p1_ca_w_0_140_s_0_210 = 3.12e-05  mcm2p1_cc_w_0_140_s_0_210 = 1.11e-10  mcm2p1_cf_w_0_140_s_0_210 = 2.93e-12
+ mcm2p1_ca_w_0_140_s_0_280 = 3.12e-05  mcm2p1_cc_w_0_140_s_0_280 = 9.50e-11  mcm2p1_cf_w_0_140_s_0_280 = 3.99e-12
+ mcm2p1_ca_w_0_140_s_0_350 = 3.12e-05  mcm2p1_cc_w_0_140_s_0_350 = 8.21e-11  mcm2p1_cf_w_0_140_s_0_350 = 5.03e-12
+ mcm2p1_ca_w_0_140_s_0_420 = 3.12e-05  mcm2p1_cc_w_0_140_s_0_420 = 7.16e-11  mcm2p1_cf_w_0_140_s_0_420 = 6.09e-12
+ mcm2p1_ca_w_0_140_s_0_560 = 3.12e-05  mcm2p1_cc_w_0_140_s_0_560 = 5.67e-11  mcm2p1_cf_w_0_140_s_0_560 = 8.03e-12
+ mcm2p1_ca_w_0_140_s_0_840 = 3.12e-05  mcm2p1_cc_w_0_140_s_0_840 = 4.08e-11  mcm2p1_cf_w_0_140_s_0_840 = 1.16e-11
+ mcm2p1_ca_w_0_140_s_1_540 = 3.12e-05  mcm2p1_cc_w_0_140_s_1_540 = 2.37e-11  mcm2p1_cf_w_0_140_s_1_540 = 1.91e-11
+ mcm2p1_ca_w_0_140_s_3_500 = 3.12e-05  mcm2p1_cc_w_0_140_s_3_500 = 9.08e-12  mcm2p1_cf_w_0_140_s_3_500 = 3.03e-11
+ mcm2p1_ca_w_1_120_s_0_140 = 3.12e-05  mcm2p1_cc_w_1_120_s_0_140 = 1.46e-10  mcm2p1_cf_w_1_120_s_0_140 = 1.92e-12
+ mcm2p1_ca_w_1_120_s_0_175 = 3.12e-05  mcm2p1_cc_w_1_120_s_0_175 = 1.39e-10  mcm2p1_cf_w_1_120_s_0_175 = 2.47e-12
+ mcm2p1_ca_w_1_120_s_0_210 = 3.12e-05  mcm2p1_cc_w_1_120_s_0_210 = 1.32e-10  mcm2p1_cf_w_1_120_s_0_210 = 3.01e-12
+ mcm2p1_ca_w_1_120_s_0_280 = 3.12e-05  mcm2p1_cc_w_1_120_s_0_280 = 1.14e-10  mcm2p1_cf_w_1_120_s_0_280 = 4.06e-12
+ mcm2p1_ca_w_1_120_s_0_350 = 3.12e-05  mcm2p1_cc_w_1_120_s_0_350 = 9.87e-11  mcm2p1_cf_w_1_120_s_0_350 = 5.10e-12
+ mcm2p1_ca_w_1_120_s_0_420 = 3.12e-05  mcm2p1_cc_w_1_120_s_0_420 = 8.69e-11  mcm2p1_cf_w_1_120_s_0_420 = 6.13e-12
+ mcm2p1_ca_w_1_120_s_0_560 = 3.12e-05  mcm2p1_cc_w_1_120_s_0_560 = 6.98e-11  mcm2p1_cf_w_1_120_s_0_560 = 8.12e-12
+ mcm2p1_ca_w_1_120_s_0_840 = 3.12e-05  mcm2p1_cc_w_1_120_s_0_840 = 5.13e-11  mcm2p1_cf_w_1_120_s_0_840 = 1.18e-11
+ mcm2p1_ca_w_1_120_s_1_540 = 3.12e-05  mcm2p1_cc_w_1_120_s_1_540 = 3.14e-11  mcm2p1_cf_w_1_120_s_1_540 = 1.95e-11
+ mcm2p1_ca_w_1_120_s_3_500 = 3.12e-05  mcm2p1_cc_w_1_120_s_3_500 = 1.35e-11  mcm2p1_cf_w_1_120_s_3_500 = 3.22e-11
+ mcm2l1_ca_w_0_140_s_0_140 = 4.60e-05  mcm2l1_cc_w_0_140_s_0_140 = 1.20e-10  mcm2l1_cf_w_0_140_s_0_140 = 2.67e-12
+ mcm2l1_ca_w_0_140_s_0_175 = 4.60e-05  mcm2l1_cc_w_0_140_s_0_175 = 1.14e-10  mcm2l1_cf_w_0_140_s_0_175 = 3.47e-12
+ mcm2l1_ca_w_0_140_s_0_210 = 4.60e-05  mcm2l1_cc_w_0_140_s_0_210 = 1.09e-10  mcm2l1_cf_w_0_140_s_0_210 = 4.26e-12
+ mcm2l1_ca_w_0_140_s_0_280 = 4.60e-05  mcm2l1_cc_w_0_140_s_0_280 = 9.39e-11  mcm2l1_cf_w_0_140_s_0_280 = 5.81e-12
+ mcm2l1_ca_w_0_140_s_0_350 = 4.60e-05  mcm2l1_cc_w_0_140_s_0_350 = 7.97e-11  mcm2l1_cf_w_0_140_s_0_350 = 7.31e-12
+ mcm2l1_ca_w_0_140_s_0_420 = 4.60e-05  mcm2l1_cc_w_0_140_s_0_420 = 6.87e-11  mcm2l1_cf_w_0_140_s_0_420 = 8.82e-12
+ mcm2l1_ca_w_0_140_s_0_560 = 4.60e-05  mcm2l1_cc_w_0_140_s_0_560 = 5.36e-11  mcm2l1_cf_w_0_140_s_0_560 = 1.15e-11
+ mcm2l1_ca_w_0_140_s_0_840 = 4.60e-05  mcm2l1_cc_w_0_140_s_0_840 = 3.74e-11  mcm2l1_cf_w_0_140_s_0_840 = 1.65e-11
+ mcm2l1_ca_w_0_140_s_1_540 = 4.60e-05  mcm2l1_cc_w_0_140_s_1_540 = 2.03e-11  mcm2l1_cf_w_0_140_s_1_540 = 2.58e-11
+ mcm2l1_ca_w_0_140_s_3_500 = 4.60e-05  mcm2l1_cc_w_0_140_s_3_500 = 6.86e-12  mcm2l1_cf_w_0_140_s_3_500 = 3.71e-11
+ mcm2l1_ca_w_1_120_s_0_140 = 4.60e-05  mcm2l1_cc_w_1_120_s_0_140 = 1.42e-10  mcm2l1_cf_w_1_120_s_0_140 = 2.71e-12
+ mcm2l1_ca_w_1_120_s_0_175 = 4.60e-05  mcm2l1_cc_w_1_120_s_0_175 = 1.35e-10  mcm2l1_cf_w_1_120_s_0_175 = 3.51e-12
+ mcm2l1_ca_w_1_120_s_0_210 = 4.60e-05  mcm2l1_cc_w_1_120_s_0_210 = 1.27e-10  mcm2l1_cf_w_1_120_s_0_210 = 4.29e-12
+ mcm2l1_ca_w_1_120_s_0_280 = 4.60e-05  mcm2l1_cc_w_1_120_s_0_280 = 1.10e-10  mcm2l1_cf_w_1_120_s_0_280 = 5.84e-12
+ mcm2l1_ca_w_1_120_s_0_350 = 4.60e-05  mcm2l1_cc_w_1_120_s_0_350 = 9.48e-11  mcm2l1_cf_w_1_120_s_0_350 = 7.35e-12
+ mcm2l1_ca_w_1_120_s_0_420 = 4.60e-05  mcm2l1_cc_w_1_120_s_0_420 = 8.26e-11  mcm2l1_cf_w_1_120_s_0_420 = 8.81e-12
+ mcm2l1_ca_w_1_120_s_0_560 = 4.60e-05  mcm2l1_cc_w_1_120_s_0_560 = 6.56e-11  mcm2l1_cf_w_1_120_s_0_560 = 1.16e-11
+ mcm2l1_ca_w_1_120_s_0_840 = 4.60e-05  mcm2l1_cc_w_1_120_s_0_840 = 4.72e-11  mcm2l1_cf_w_1_120_s_0_840 = 1.66e-11
+ mcm2l1_ca_w_1_120_s_1_540 = 4.60e-05  mcm2l1_cc_w_1_120_s_1_540 = 2.76e-11  mcm2l1_cf_w_1_120_s_1_540 = 2.62e-11
+ mcm2l1_ca_w_1_120_s_3_500 = 4.60e-05  mcm2l1_cc_w_1_120_s_3_500 = 1.10e-11  mcm2l1_cf_w_1_120_s_3_500 = 3.94e-11
+ mcm2m1_ca_w_0_140_s_0_140 = 2.18e-04  mcm2m1_cc_w_0_140_s_0_140 = 1.08e-10  mcm2m1_cf_w_0_140_s_0_140 = 1.14e-11
+ mcm2m1_ca_w_0_140_s_0_175 = 2.18e-04  mcm2m1_cc_w_0_140_s_0_175 = 1.01e-10  mcm2m1_cf_w_0_140_s_0_175 = 1.52e-11
+ mcm2m1_ca_w_0_140_s_0_210 = 2.18e-04  mcm2m1_cc_w_0_140_s_0_210 = 9.47e-11  mcm2m1_cf_w_0_140_s_0_210 = 1.87e-11
+ mcm2m1_ca_w_0_140_s_0_280 = 2.18e-04  mcm2m1_cc_w_0_140_s_0_280 = 7.92e-11  mcm2m1_cf_w_0_140_s_0_280 = 2.50e-11
+ mcm2m1_ca_w_0_140_s_0_350 = 2.18e-04  mcm2m1_cc_w_0_140_s_0_350 = 6.51e-11  mcm2m1_cf_w_0_140_s_0_350 = 3.05e-11
+ mcm2m1_ca_w_0_140_s_0_420 = 2.18e-04  mcm2m1_cc_w_0_140_s_0_420 = 5.39e-11  mcm2m1_cf_w_0_140_s_0_420 = 3.53e-11
+ mcm2m1_ca_w_0_140_s_0_560 = 2.18e-04  mcm2m1_cc_w_0_140_s_0_560 = 3.92e-11  mcm2m1_cf_w_0_140_s_0_560 = 4.30e-11
+ mcm2m1_ca_w_0_140_s_0_840 = 2.18e-04  mcm2m1_cc_w_0_140_s_0_840 = 2.45e-11  mcm2m1_cf_w_0_140_s_0_840 = 5.35e-11
+ mcm2m1_ca_w_0_140_s_1_540 = 2.18e-04  mcm2m1_cc_w_0_140_s_1_540 = 1.06e-11  mcm2m1_cf_w_0_140_s_1_540 = 6.60e-11
+ mcm2m1_ca_w_0_140_s_3_500 = 2.18e-04  mcm2m1_cc_w_0_140_s_3_500 = 2.90e-12  mcm2m1_cf_w_0_140_s_3_500 = 7.43e-11
+ mcm2m1_ca_w_1_120_s_0_140 = 2.18e-04  mcm2m1_cc_w_1_120_s_0_140 = 1.25e-10  mcm2m1_cf_w_1_120_s_0_140 = 1.14e-11
+ mcm2m1_ca_w_1_120_s_0_175 = 2.18e-04  mcm2m1_cc_w_1_120_s_0_175 = 1.18e-10  mcm2m1_cf_w_1_120_s_0_175 = 1.52e-11
+ mcm2m1_ca_w_1_120_s_0_210 = 2.18e-04  mcm2m1_cc_w_1_120_s_0_210 = 1.10e-10  mcm2m1_cf_w_1_120_s_0_210 = 1.87e-11
+ mcm2m1_ca_w_1_120_s_0_280 = 2.18e-04  mcm2m1_cc_w_1_120_s_0_280 = 9.29e-11  mcm2m1_cf_w_1_120_s_0_280 = 2.50e-11
+ mcm2m1_ca_w_1_120_s_0_350 = 2.18e-04  mcm2m1_cc_w_1_120_s_0_350 = 7.84e-11  mcm2m1_cf_w_1_120_s_0_350 = 3.05e-11
+ mcm2m1_ca_w_1_120_s_0_420 = 2.18e-04  mcm2m1_cc_w_1_120_s_0_420 = 6.65e-11  mcm2m1_cf_w_1_120_s_0_420 = 3.53e-11
+ mcm2m1_ca_w_1_120_s_0_560 = 2.18e-04  mcm2m1_cc_w_1_120_s_0_560 = 5.05e-11  mcm2m1_cf_w_1_120_s_0_560 = 4.30e-11
+ mcm2m1_ca_w_1_120_s_0_840 = 2.18e-04  mcm2m1_cc_w_1_120_s_0_840 = 3.38e-11  mcm2m1_cf_w_1_120_s_0_840 = 5.36e-11
+ mcm2m1_ca_w_1_120_s_1_540 = 2.18e-04  mcm2m1_cc_w_1_120_s_1_540 = 1.77e-11  mcm2m1_cf_w_1_120_s_1_540 = 6.73e-11
+ mcm2m1_ca_w_1_120_s_3_500 = 2.18e-04  mcm2m1_cc_w_1_120_s_3_500 = 6.20e-12  mcm2m1_cf_w_1_120_s_3_500 = 7.89e-11
+ mcm3f_ca_w_0_300_s_0_300 = 1.49e-05  mcm3f_cc_w_0_300_s_0_300 = 1.18e-10  mcm3f_cf_w_0_300_s_0_300 = 1.96e-12
+ mcm3f_ca_w_0_300_s_0_360 = 1.49e-05  mcm3f_cc_w_0_300_s_0_360 = 1.10e-10  mcm3f_cf_w_0_300_s_0_360 = 2.40e-12
+ mcm3f_ca_w_0_300_s_0_450 = 1.49e-05  mcm3f_cc_w_0_300_s_0_450 = 9.84e-11  mcm3f_cf_w_0_300_s_0_450 = 3.06e-12
+ mcm3f_ca_w_0_300_s_0_600 = 1.49e-05  mcm3f_cc_w_0_300_s_0_600 = 8.33e-11  mcm3f_cf_w_0_300_s_0_600 = 4.13e-12
+ mcm3f_ca_w_0_300_s_0_800 = 1.49e-05  mcm3f_cc_w_0_300_s_0_800 = 6.94e-11  mcm3f_cf_w_0_300_s_0_800 = 5.44e-12
+ mcm3f_ca_w_0_300_s_1_000 = 1.49e-05  mcm3f_cc_w_0_300_s_1_000 = 5.94e-11  mcm3f_cf_w_0_300_s_1_000 = 6.76e-12
+ mcm3f_ca_w_0_300_s_1_200 = 1.49e-05  mcm3f_cc_w_0_300_s_1_200 = 5.16e-11  mcm3f_cf_w_0_300_s_1_200 = 8.03e-12
+ mcm3f_ca_w_0_300_s_2_100 = 1.49e-05  mcm3f_cc_w_0_300_s_2_100 = 3.31e-11  mcm3f_cf_w_0_300_s_2_100 = 1.35e-11
+ mcm3f_ca_w_0_300_s_3_300 = 1.49e-05  mcm3f_cc_w_0_300_s_3_300 = 2.26e-11  mcm3f_cf_w_0_300_s_3_300 = 1.87e-11
+ mcm3f_ca_w_0_300_s_9_000 = 1.49e-05  mcm3f_cc_w_0_300_s_9_000 = 6.59e-12  mcm3f_cf_w_0_300_s_9_000 = 3.11e-11
+ mcm3f_ca_w_2_400_s_0_300 = 1.49e-05  mcm3f_cc_w_2_400_s_0_300 = 1.43e-10  mcm3f_cf_w_2_400_s_0_300 = 2.01e-12
+ mcm3f_ca_w_2_400_s_0_360 = 1.49e-05  mcm3f_cc_w_2_400_s_0_360 = 1.33e-10  mcm3f_cf_w_2_400_s_0_360 = 2.44e-12
+ mcm3f_ca_w_2_400_s_0_450 = 1.49e-05  mcm3f_cc_w_2_400_s_0_450 = 1.20e-10  mcm3f_cf_w_2_400_s_0_450 = 3.09e-12
+ mcm3f_ca_w_2_400_s_0_600 = 1.49e-05  mcm3f_cc_w_2_400_s_0_600 = 1.02e-10  mcm3f_cf_w_2_400_s_0_600 = 4.14e-12
+ mcm3f_ca_w_2_400_s_0_800 = 1.49e-05  mcm3f_cc_w_2_400_s_0_800 = 8.64e-11  mcm3f_cf_w_2_400_s_0_800 = 5.51e-12
+ mcm3f_ca_w_2_400_s_1_000 = 1.49e-05  mcm3f_cc_w_2_400_s_1_000 = 7.44e-11  mcm3f_cf_w_2_400_s_1_000 = 6.85e-12
+ mcm3f_ca_w_2_400_s_1_200 = 1.49e-05  mcm3f_cc_w_2_400_s_1_200 = 6.57e-11  mcm3f_cf_w_2_400_s_1_200 = 8.13e-12
+ mcm3f_ca_w_2_400_s_2_100 = 1.49e-05  mcm3f_cc_w_2_400_s_2_100 = 4.40e-11  mcm3f_cf_w_2_400_s_2_100 = 1.34e-11
+ mcm3f_ca_w_2_400_s_3_300 = 1.49e-05  mcm3f_cc_w_2_400_s_3_300 = 3.08e-11  mcm3f_cf_w_2_400_s_3_300 = 1.92e-11
+ mcm3f_ca_w_2_400_s_9_000 = 1.49e-05  mcm3f_cc_w_2_400_s_9_000 = 1.04e-11  mcm3f_cf_w_2_400_s_9_000 = 3.39e-11
+ mcm3d_ca_w_0_300_s_0_300 = 1.67e-05  mcm3d_cc_w_0_300_s_0_300 = 1.18e-10  mcm3d_cf_w_0_300_s_0_300 = 2.19e-12
+ mcm3d_ca_w_0_300_s_0_360 = 1.67e-05  mcm3d_cc_w_0_300_s_0_360 = 1.10e-10  mcm3d_cf_w_0_300_s_0_360 = 2.67e-12
+ mcm3d_ca_w_0_300_s_0_450 = 1.67e-05  mcm3d_cc_w_0_300_s_0_450 = 9.79e-11  mcm3d_cf_w_0_300_s_0_450 = 3.40e-12
+ mcm3d_ca_w_0_300_s_0_600 = 1.67e-05  mcm3d_cc_w_0_300_s_0_600 = 8.28e-11  mcm3d_cf_w_0_300_s_0_600 = 4.59e-12
+ mcm3d_ca_w_0_300_s_0_800 = 1.67e-05  mcm3d_cc_w_0_300_s_0_800 = 6.87e-11  mcm3d_cf_w_0_300_s_0_800 = 6.03e-12
+ mcm3d_ca_w_0_300_s_1_000 = 1.67e-05  mcm3d_cc_w_0_300_s_1_000 = 5.85e-11  mcm3d_cf_w_0_300_s_1_000 = 7.46e-12
+ mcm3d_ca_w_0_300_s_1_200 = 1.67e-05  mcm3d_cc_w_0_300_s_1_200 = 5.08e-11  mcm3d_cf_w_0_300_s_1_200 = 8.87e-12
+ mcm3d_ca_w_0_300_s_2_100 = 1.67e-05  mcm3d_cc_w_0_300_s_2_100 = 3.22e-11  mcm3d_cf_w_0_300_s_2_100 = 1.48e-11
+ mcm3d_ca_w_0_300_s_3_300 = 1.67e-05  mcm3d_cc_w_0_300_s_3_300 = 2.17e-11  mcm3d_cf_w_0_300_s_3_300 = 2.03e-11
+ mcm3d_ca_w_0_300_s_9_000 = 1.67e-05  mcm3d_cc_w_0_300_s_9_000 = 6.05e-12  mcm3d_cf_w_0_300_s_9_000 = 3.27e-11
+ mcm3d_ca_w_2_400_s_0_300 = 1.67e-05  mcm3d_cc_w_2_400_s_0_300 = 1.42e-10  mcm3d_cf_w_2_400_s_0_300 = 2.24e-12
+ mcm3d_ca_w_2_400_s_0_360 = 1.67e-05  mcm3d_cc_w_2_400_s_0_360 = 1.32e-10  mcm3d_cf_w_2_400_s_0_360 = 2.72e-12
+ mcm3d_ca_w_2_400_s_0_450 = 1.67e-05  mcm3d_cc_w_2_400_s_0_450 = 1.19e-10  mcm3d_cf_w_2_400_s_0_450 = 3.44e-12
+ mcm3d_ca_w_2_400_s_0_600 = 1.67e-05  mcm3d_cc_w_2_400_s_0_600 = 1.01e-10  mcm3d_cf_w_2_400_s_0_600 = 4.60e-12
+ mcm3d_ca_w_2_400_s_0_800 = 1.67e-05  mcm3d_cc_w_2_400_s_0_800 = 8.52e-11  mcm3d_cf_w_2_400_s_0_800 = 6.11e-12
+ mcm3d_ca_w_2_400_s_1_000 = 1.67e-05  mcm3d_cc_w_2_400_s_1_000 = 7.33e-11  mcm3d_cf_w_2_400_s_1_000 = 7.59e-12
+ mcm3d_ca_w_2_400_s_1_200 = 1.67e-05  mcm3d_cc_w_2_400_s_1_200 = 6.44e-11  mcm3d_cf_w_2_400_s_1_200 = 9.00e-12
+ mcm3d_ca_w_2_400_s_2_100 = 1.67e-05  mcm3d_cc_w_2_400_s_2_100 = 4.28e-11  mcm3d_cf_w_2_400_s_2_100 = 1.47e-11
+ mcm3d_ca_w_2_400_s_3_300 = 1.67e-05  mcm3d_cc_w_2_400_s_3_300 = 2.97e-11  mcm3d_cf_w_2_400_s_3_300 = 2.09e-11
+ mcm3d_ca_w_2_400_s_9_000 = 1.67e-05  mcm3d_cc_w_2_400_s_9_000 = 9.75e-12  mcm3d_cf_w_2_400_s_9_000 = 3.57e-11
+ mcm3p1_ca_w_0_300_s_0_300 = 1.92e-05  mcm3p1_cc_w_0_300_s_0_300 = 1.17e-10  mcm3p1_cf_w_0_300_s_0_300 = 2.53e-12
+ mcm3p1_ca_w_0_300_s_0_360 = 1.92e-05  mcm3p1_cc_w_0_300_s_0_360 = 1.09e-10  mcm3p1_cf_w_0_300_s_0_360 = 3.08e-12
+ mcm3p1_ca_w_0_300_s_0_450 = 1.92e-05  mcm3p1_cc_w_0_300_s_0_450 = 9.72e-11  mcm3p1_cf_w_0_300_s_0_450 = 3.91e-12
+ mcm3p1_ca_w_0_300_s_0_600 = 1.92e-05  mcm3p1_cc_w_0_300_s_0_600 = 8.19e-11  mcm3p1_cf_w_0_300_s_0_600 = 5.26e-12
+ mcm3p1_ca_w_0_300_s_0_800 = 1.92e-05  mcm3p1_cc_w_0_300_s_0_800 = 6.79e-11  mcm3p1_cf_w_0_300_s_0_800 = 6.92e-12
+ mcm3p1_ca_w_0_300_s_1_000 = 1.92e-05  mcm3p1_cc_w_0_300_s_1_000 = 5.74e-11  mcm3p1_cf_w_0_300_s_1_000 = 8.55e-12
+ mcm3p1_ca_w_0_300_s_1_200 = 1.92e-05  mcm3p1_cc_w_0_300_s_1_200 = 4.97e-11  mcm3p1_cf_w_0_300_s_1_200 = 1.01e-11
+ mcm3p1_ca_w_0_300_s_2_100 = 1.92e-05  mcm3p1_cc_w_0_300_s_2_100 = 3.09e-11  mcm3p1_cf_w_0_300_s_2_100 = 1.67e-11
+ mcm3p1_ca_w_0_300_s_3_300 = 1.92e-05  mcm3p1_cc_w_0_300_s_3_300 = 2.04e-11  mcm3p1_cf_w_0_300_s_3_300 = 2.26e-11
+ mcm3p1_ca_w_0_300_s_9_000 = 1.92e-05  mcm3p1_cc_w_0_300_s_9_000 = 5.45e-12  mcm3p1_cf_w_0_300_s_9_000 = 3.48e-11
+ mcm3p1_ca_w_2_400_s_0_300 = 1.92e-05  mcm3p1_cc_w_2_400_s_0_300 = 1.40e-10  mcm3p1_cf_w_2_400_s_0_300 = 2.62e-12
+ mcm3p1_ca_w_2_400_s_0_360 = 1.92e-05  mcm3p1_cc_w_2_400_s_0_360 = 1.30e-10  mcm3p1_cf_w_2_400_s_0_360 = 3.16e-12
+ mcm3p1_ca_w_2_400_s_0_450 = 1.92e-05  mcm3p1_cc_w_2_400_s_0_450 = 1.17e-10  mcm3p1_cf_w_2_400_s_0_450 = 3.98e-12
+ mcm3p1_ca_w_2_400_s_0_600 = 1.92e-05  mcm3p1_cc_w_2_400_s_0_600 = 9.96e-11  mcm3p1_cf_w_2_400_s_0_600 = 5.31e-12
+ mcm3p1_ca_w_2_400_s_0_800 = 1.92e-05  mcm3p1_cc_w_2_400_s_0_800 = 8.37e-11  mcm3p1_cf_w_2_400_s_0_800 = 7.03e-12
+ mcm3p1_ca_w_2_400_s_1_000 = 1.92e-05  mcm3p1_cc_w_2_400_s_1_000 = 7.17e-11  mcm3p1_cf_w_2_400_s_1_000 = 8.72e-12
+ mcm3p1_ca_w_2_400_s_1_200 = 1.92e-05  mcm3p1_cc_w_2_400_s_1_200 = 6.30e-11  mcm3p1_cf_w_2_400_s_1_200 = 1.03e-11
+ mcm3p1_ca_w_2_400_s_2_100 = 1.92e-05  mcm3p1_cc_w_2_400_s_2_100 = 4.13e-11  mcm3p1_cf_w_2_400_s_2_100 = 1.66e-11
+ mcm3p1_ca_w_2_400_s_3_300 = 1.92e-05  mcm3p1_cc_w_2_400_s_3_300 = 2.82e-11  mcm3p1_cf_w_2_400_s_3_300 = 2.32e-11
+ mcm3p1_ca_w_2_400_s_9_000 = 1.92e-05  mcm3p1_cc_w_2_400_s_9_000 = 9.00e-12  mcm3p1_cf_w_2_400_s_9_000 = 3.82e-11
+ mcm3l1_ca_w_0_300_s_0_300 = 2.40e-05  mcm3l1_cc_w_0_300_s_0_300 = 1.16e-10  mcm3l1_cf_w_0_300_s_0_300 = 3.12e-12
+ mcm3l1_ca_w_0_300_s_0_360 = 2.40e-05  mcm3l1_cc_w_0_300_s_0_360 = 1.07e-10  mcm3l1_cf_w_0_300_s_0_360 = 3.79e-12
+ mcm3l1_ca_w_0_300_s_0_450 = 2.40e-05  mcm3l1_cc_w_0_300_s_0_450 = 9.56e-11  mcm3l1_cf_w_0_300_s_0_450 = 4.81e-12
+ mcm3l1_ca_w_0_300_s_0_600 = 2.40e-05  mcm3l1_cc_w_0_300_s_0_600 = 8.05e-11  mcm3l1_cf_w_0_300_s_0_600 = 6.45e-12
+ mcm3l1_ca_w_0_300_s_0_800 = 2.40e-05  mcm3l1_cc_w_0_300_s_0_800 = 6.63e-11  mcm3l1_cf_w_0_300_s_0_800 = 8.46e-12
+ mcm3l1_ca_w_0_300_s_1_000 = 2.40e-05  mcm3l1_cc_w_0_300_s_1_000 = 5.58e-11  mcm3l1_cf_w_0_300_s_1_000 = 1.04e-11
+ mcm3l1_ca_w_0_300_s_1_200 = 2.40e-05  mcm3l1_cc_w_0_300_s_1_200 = 4.80e-11  mcm3l1_cf_w_0_300_s_1_200 = 1.23e-11
+ mcm3l1_ca_w_0_300_s_2_100 = 2.40e-05  mcm3l1_cc_w_0_300_s_2_100 = 2.90e-11  mcm3l1_cf_w_0_300_s_2_100 = 1.98e-11
+ mcm3l1_ca_w_0_300_s_3_300 = 2.40e-05  mcm3l1_cc_w_0_300_s_3_300 = 1.86e-11  mcm3l1_cf_w_0_300_s_3_300 = 2.61e-11
+ mcm3l1_ca_w_0_300_s_9_000 = 2.40e-05  mcm3l1_cc_w_0_300_s_9_000 = 4.63e-12  mcm3l1_cf_w_0_300_s_9_000 = 3.80e-11
+ mcm3l1_ca_w_2_400_s_0_300 = 2.40e-05  mcm3l1_cc_w_2_400_s_0_300 = 1.38e-10  mcm3l1_cf_w_2_400_s_0_300 = 3.16e-12
+ mcm3l1_ca_w_2_400_s_0_360 = 2.40e-05  mcm3l1_cc_w_2_400_s_0_360 = 1.28e-10  mcm3l1_cf_w_2_400_s_0_360 = 3.84e-12
+ mcm3l1_ca_w_2_400_s_0_450 = 2.40e-05  mcm3l1_cc_w_2_400_s_0_450 = 1.14e-10  mcm3l1_cf_w_2_400_s_0_450 = 4.84e-12
+ mcm3l1_ca_w_2_400_s_0_600 = 2.40e-05  mcm3l1_cc_w_2_400_s_0_600 = 9.72e-11  mcm3l1_cf_w_2_400_s_0_600 = 6.46e-12
+ mcm3l1_ca_w_2_400_s_0_800 = 2.40e-05  mcm3l1_cc_w_2_400_s_0_800 = 8.14e-11  mcm3l1_cf_w_2_400_s_0_800 = 8.53e-12
+ mcm3l1_ca_w_2_400_s_1_000 = 2.40e-05  mcm3l1_cc_w_2_400_s_1_000 = 6.92e-11  mcm3l1_cf_w_2_400_s_1_000 = 1.05e-11
+ mcm3l1_ca_w_2_400_s_1_200 = 2.40e-05  mcm3l1_cc_w_2_400_s_1_200 = 6.05e-11  mcm3l1_cf_w_2_400_s_1_200 = 1.24e-11
+ mcm3l1_ca_w_2_400_s_2_100 = 2.40e-05  mcm3l1_cc_w_2_400_s_2_100 = 3.92e-11  mcm3l1_cf_w_2_400_s_2_100 = 1.97e-11
+ mcm3l1_ca_w_2_400_s_3_300 = 2.40e-05  mcm3l1_cc_w_2_400_s_3_300 = 2.62e-11  mcm3l1_cf_w_2_400_s_3_300 = 2.69e-11
+ mcm3l1_ca_w_2_400_s_9_000 = 2.40e-05  mcm3l1_cc_w_2_400_s_9_000 = 7.95e-12  mcm3l1_cf_w_2_400_s_9_000 = 4.17e-11
+ mcm3m1_ca_w_0_300_s_0_300 = 4.08e-05  mcm3m1_cc_w_0_300_s_0_300 = 1.13e-10  mcm3m1_cf_w_0_300_s_0_300 = 5.19e-12
+ mcm3m1_ca_w_0_300_s_0_360 = 4.08e-05  mcm3m1_cc_w_0_300_s_0_360 = 1.03e-10  mcm3m1_cf_w_0_300_s_0_360 = 6.29e-12
+ mcm3m1_ca_w_0_300_s_0_450 = 4.08e-05  mcm3m1_cc_w_0_300_s_0_450 = 9.16e-11  mcm3m1_cf_w_0_300_s_0_450 = 7.90e-12
+ mcm3m1_ca_w_0_300_s_0_600 = 4.08e-05  mcm3m1_cc_w_0_300_s_0_600 = 7.63e-11  mcm3m1_cf_w_0_300_s_0_600 = 1.05e-11
+ mcm3m1_ca_w_0_300_s_0_800 = 4.08e-05  mcm3m1_cc_w_0_300_s_0_800 = 6.18e-11  mcm3m1_cf_w_0_300_s_0_800 = 1.36e-11
+ mcm3m1_ca_w_0_300_s_1_000 = 4.08e-05  mcm3m1_cc_w_0_300_s_1_000 = 5.10e-11  mcm3m1_cf_w_0_300_s_1_000 = 1.64e-11
+ mcm3m1_ca_w_0_300_s_1_200 = 4.08e-05  mcm3m1_cc_w_0_300_s_1_200 = 4.32e-11  mcm3m1_cf_w_0_300_s_1_200 = 1.91e-11
+ mcm3m1_ca_w_0_300_s_2_100 = 4.08e-05  mcm3m1_cc_w_0_300_s_2_100 = 2.43e-11  mcm3m1_cf_w_0_300_s_2_100 = 2.88e-11
+ mcm3m1_ca_w_0_300_s_3_300 = 4.08e-05  mcm3m1_cc_w_0_300_s_3_300 = 1.47e-11  mcm3m1_cf_w_0_300_s_3_300 = 3.58e-11
+ mcm3m1_ca_w_0_300_s_9_000 = 4.08e-05  mcm3m1_cc_w_0_300_s_9_000 = 3.25e-12  mcm3m1_cf_w_0_300_s_9_000 = 4.63e-11
+ mcm3m1_ca_w_2_400_s_0_300 = 4.08e-05  mcm3m1_cc_w_2_400_s_0_300 = 1.32e-10  mcm3m1_cf_w_2_400_s_0_300 = 5.19e-12
+ mcm3m1_ca_w_2_400_s_0_360 = 4.08e-05  mcm3m1_cc_w_2_400_s_0_360 = 1.22e-10  mcm3m1_cf_w_2_400_s_0_360 = 6.29e-12
+ mcm3m1_ca_w_2_400_s_0_450 = 4.08e-05  mcm3m1_cc_w_2_400_s_0_450 = 1.09e-10  mcm3m1_cf_w_2_400_s_0_450 = 7.90e-12
+ mcm3m1_ca_w_2_400_s_0_600 = 4.08e-05  mcm3m1_cc_w_2_400_s_0_600 = 9.16e-11  mcm3m1_cf_w_2_400_s_0_600 = 1.05e-11
+ mcm3m1_ca_w_2_400_s_0_800 = 4.08e-05  mcm3m1_cc_w_2_400_s_0_800 = 7.57e-11  mcm3m1_cf_w_2_400_s_0_800 = 1.36e-11
+ mcm3m1_ca_w_2_400_s_1_000 = 4.08e-05  mcm3m1_cc_w_2_400_s_1_000 = 6.38e-11  mcm3m1_cf_w_2_400_s_1_000 = 1.65e-11
+ mcm3m1_ca_w_2_400_s_1_200 = 4.08e-05  mcm3m1_cc_w_2_400_s_1_200 = 5.51e-11  mcm3m1_cf_w_2_400_s_1_200 = 1.91e-11
+ mcm3m1_ca_w_2_400_s_2_100 = 4.08e-05  mcm3m1_cc_w_2_400_s_2_100 = 3.43e-11  mcm3m1_cf_w_2_400_s_2_100 = 2.86e-11
+ mcm3m1_ca_w_2_400_s_3_300 = 4.08e-05  mcm3m1_cc_w_2_400_s_3_300 = 2.22e-11  mcm3m1_cf_w_2_400_s_3_300 = 3.68e-11
+ mcm3m1_ca_w_2_400_s_9_000 = 4.08e-05  mcm3m1_cc_w_2_400_s_9_000 = 6.15e-12  mcm3m1_cf_w_2_400_s_9_000 = 5.08e-11
+ mcm3m2_ca_w_0_300_s_0_300 = 1.12e-04  mcm3m2_cc_w_0_300_s_0_300 = 1.03e-10  mcm3m2_cf_w_0_300_s_0_300 = 1.32e-11
+ mcm3m2_ca_w_0_300_s_0_360 = 1.12e-04  mcm3m2_cc_w_0_300_s_0_360 = 9.37e-11  mcm3m2_cf_w_0_300_s_0_360 = 1.57e-11
+ mcm3m2_ca_w_0_300_s_0_450 = 1.12e-04  mcm3m2_cc_w_0_300_s_0_450 = 8.21e-11  mcm3m2_cf_w_0_300_s_0_450 = 1.91e-11
+ mcm3m2_ca_w_0_300_s_0_600 = 1.12e-04  mcm3m2_cc_w_0_300_s_0_600 = 6.66e-11  mcm3m2_cf_w_0_300_s_0_600 = 2.42e-11
+ mcm3m2_ca_w_0_300_s_0_800 = 1.12e-04  mcm3m2_cc_w_0_300_s_0_800 = 5.27e-11  mcm3m2_cf_w_0_300_s_0_800 = 2.96e-11
+ mcm3m2_ca_w_0_300_s_1_000 = 1.12e-04  mcm3m2_cc_w_0_300_s_1_000 = 4.25e-11  mcm3m2_cf_w_0_300_s_1_000 = 3.42e-11
+ mcm3m2_ca_w_0_300_s_1_200 = 1.12e-04  mcm3m2_cc_w_0_300_s_1_200 = 3.51e-11  mcm3m2_cf_w_0_300_s_1_200 = 3.80e-11
+ mcm3m2_ca_w_0_300_s_2_100 = 1.12e-04  mcm3m2_cc_w_0_300_s_2_100 = 1.78e-11  mcm3m2_cf_w_0_300_s_2_100 = 4.98e-11
+ mcm3m2_ca_w_0_300_s_3_300 = 1.12e-04  mcm3m2_cc_w_0_300_s_3_300 = 1.01e-11  mcm3m2_cf_w_0_300_s_3_300 = 5.64e-11
+ mcm3m2_ca_w_0_300_s_9_000 = 1.12e-04  mcm3m2_cc_w_0_300_s_9_000 = 2.10e-12  mcm3m2_cf_w_0_300_s_9_000 = 6.42e-11
+ mcm3m2_ca_w_2_400_s_0_300 = 1.12e-04  mcm3m2_cc_w_2_400_s_0_300 = 1.21e-10  mcm3m2_cf_w_2_400_s_0_300 = 1.32e-11
+ mcm3m2_ca_w_2_400_s_0_360 = 1.12e-04  mcm3m2_cc_w_2_400_s_0_360 = 1.11e-10  mcm3m2_cf_w_2_400_s_0_360 = 1.57e-11
+ mcm3m2_ca_w_2_400_s_0_450 = 1.12e-04  mcm3m2_cc_w_2_400_s_0_450 = 9.80e-11  mcm3m2_cf_w_2_400_s_0_450 = 1.91e-11
+ mcm3m2_ca_w_2_400_s_0_600 = 1.12e-04  mcm3m2_cc_w_2_400_s_0_600 = 8.16e-11  mcm3m2_cf_w_2_400_s_0_600 = 2.41e-11
+ mcm3m2_ca_w_2_400_s_0_800 = 1.12e-04  mcm3m2_cc_w_2_400_s_0_800 = 6.61e-11  mcm3m2_cf_w_2_400_s_0_800 = 2.96e-11
+ mcm3m2_ca_w_2_400_s_1_000 = 1.12e-04  mcm3m2_cc_w_2_400_s_1_000 = 5.49e-11  mcm3m2_cf_w_2_400_s_1_000 = 3.42e-11
+ mcm3m2_ca_w_2_400_s_1_200 = 1.12e-04  mcm3m2_cc_w_2_400_s_1_200 = 4.68e-11  mcm3m2_cf_w_2_400_s_1_200 = 3.79e-11
+ mcm3m2_ca_w_2_400_s_2_100 = 1.12e-04  mcm3m2_cc_w_2_400_s_2_100 = 2.79e-11  mcm3m2_cf_w_2_400_s_2_100 = 4.96e-11
+ mcm3m2_ca_w_2_400_s_3_300 = 1.12e-04  mcm3m2_cc_w_2_400_s_3_300 = 1.74e-11  mcm3m2_cf_w_2_400_s_3_300 = 5.81e-11
+ mcm3m2_ca_w_2_400_s_9_000 = 1.12e-04  mcm3m2_cc_w_2_400_s_9_000 = 4.60e-12  mcm3m2_cf_w_2_400_s_9_000 = 7.02e-11
+ mcm4f_ca_w_0_300_s_0_300 = 9.99e-06  mcm4f_cc_w_0_300_s_0_300 = 1.21e-10  mcm4f_cf_w_0_300_s_0_300 = 1.32e-12
+ mcm4f_ca_w_0_300_s_0_360 = 9.99e-06  mcm4f_cc_w_0_300_s_0_360 = 1.12e-10  mcm4f_cf_w_0_300_s_0_360 = 1.61e-12
+ mcm4f_ca_w_0_300_s_0_450 = 9.99e-06  mcm4f_cc_w_0_300_s_0_450 = 1.01e-10  mcm4f_cf_w_0_300_s_0_450 = 2.07e-12
+ mcm4f_ca_w_0_300_s_0_600 = 9.99e-06  mcm4f_cc_w_0_300_s_0_600 = 8.68e-11  mcm4f_cf_w_0_300_s_0_600 = 2.81e-12
+ mcm4f_ca_w_0_300_s_0_800 = 9.99e-06  mcm4f_cc_w_0_300_s_0_800 = 7.34e-11  mcm4f_cf_w_0_300_s_0_800 = 3.70e-12
+ mcm4f_ca_w_0_300_s_1_000 = 9.99e-06  mcm4f_cc_w_0_300_s_1_000 = 6.34e-11  mcm4f_cf_w_0_300_s_1_000 = 4.61e-12
+ mcm4f_ca_w_0_300_s_1_200 = 9.99e-06  mcm4f_cc_w_0_300_s_1_200 = 5.61e-11  mcm4f_cf_w_0_300_s_1_200 = 5.51e-12
+ mcm4f_ca_w_0_300_s_2_100 = 9.99e-06  mcm4f_cc_w_0_300_s_2_100 = 3.80e-11  mcm4f_cf_w_0_300_s_2_100 = 9.53e-12
+ mcm4f_ca_w_0_300_s_3_300 = 9.99e-06  mcm4f_cc_w_0_300_s_3_300 = 2.71e-11  mcm4f_cf_w_0_300_s_3_300 = 1.36e-11
+ mcm4f_ca_w_0_300_s_9_000 = 9.99e-06  mcm4f_cc_w_0_300_s_9_000 = 9.25e-12  mcm4f_cf_w_0_300_s_9_000 = 2.55e-11
+ mcm4f_ca_w_2_400_s_0_300 = 9.99e-06  mcm4f_cc_w_2_400_s_0_300 = 1.51e-10  mcm4f_cf_w_2_400_s_0_300 = 1.35e-12
+ mcm4f_ca_w_2_400_s_0_360 = 9.99e-06  mcm4f_cc_w_2_400_s_0_360 = 1.40e-10  mcm4f_cf_w_2_400_s_0_360 = 1.64e-12
+ mcm4f_ca_w_2_400_s_0_450 = 9.99e-06  mcm4f_cc_w_2_400_s_0_450 = 1.27e-10  mcm4f_cf_w_2_400_s_0_450 = 2.07e-12
+ mcm4f_ca_w_2_400_s_0_600 = 9.99e-06  mcm4f_cc_w_2_400_s_0_600 = 1.10e-10  mcm4f_cf_w_2_400_s_0_600 = 2.79e-12
+ mcm4f_ca_w_2_400_s_0_800 = 9.99e-06  mcm4f_cc_w_2_400_s_0_800 = 9.38e-11  mcm4f_cf_w_2_400_s_0_800 = 3.73e-12
+ mcm4f_ca_w_2_400_s_1_000 = 9.99e-06  mcm4f_cc_w_2_400_s_1_000 = 8.17e-11  mcm4f_cf_w_2_400_s_1_000 = 4.67e-12
+ mcm4f_ca_w_2_400_s_1_200 = 9.99e-06  mcm4f_cc_w_2_400_s_1_200 = 7.26e-11  mcm4f_cf_w_2_400_s_1_200 = 5.57e-12
+ mcm4f_ca_w_2_400_s_2_100 = 9.99e-06  mcm4f_cc_w_2_400_s_2_100 = 5.01e-11  mcm4f_cf_w_2_400_s_2_100 = 9.40e-12
+ mcm4f_ca_w_2_400_s_3_300 = 9.99e-06  mcm4f_cc_w_2_400_s_3_300 = 3.61e-11  mcm4f_cf_w_2_400_s_3_300 = 1.39e-11
+ mcm4f_ca_w_2_400_s_9_000 = 9.99e-06  mcm4f_cc_w_2_400_s_9_000 = 1.34e-11  mcm4f_cf_w_2_400_s_9_000 = 2.76e-11
+ mcm4d_ca_w_0_300_s_0_300 = 1.07e-05  mcm4d_cc_w_0_300_s_0_300 = 1.21e-10  mcm4d_cf_w_0_300_s_0_300 = 1.41e-12
+ mcm4d_ca_w_0_300_s_0_360 = 1.07e-05  mcm4d_cc_w_0_300_s_0_360 = 1.12e-10  mcm4d_cf_w_0_300_s_0_360 = 1.73e-12
+ mcm4d_ca_w_0_300_s_0_450 = 1.07e-05  mcm4d_cc_w_0_300_s_0_450 = 1.00e-10  mcm4d_cf_w_0_300_s_0_450 = 2.22e-12
+ mcm4d_ca_w_0_300_s_0_600 = 1.07e-05  mcm4d_cc_w_0_300_s_0_600 = 8.65e-11  mcm4d_cf_w_0_300_s_0_600 = 3.01e-12
+ mcm4d_ca_w_0_300_s_0_800 = 1.07e-05  mcm4d_cc_w_0_300_s_0_800 = 7.31e-11  mcm4d_cf_w_0_300_s_0_800 = 3.96e-12
+ mcm4d_ca_w_0_300_s_1_000 = 1.07e-05  mcm4d_cc_w_0_300_s_1_000 = 6.31e-11  mcm4d_cf_w_0_300_s_1_000 = 4.94e-12
+ mcm4d_ca_w_0_300_s_1_200 = 1.07e-05  mcm4d_cc_w_0_300_s_1_200 = 5.57e-11  mcm4d_cf_w_0_300_s_1_200 = 5.90e-12
+ mcm4d_ca_w_0_300_s_2_100 = 1.07e-05  mcm4d_cc_w_0_300_s_2_100 = 3.74e-11  mcm4d_cf_w_0_300_s_2_100 = 1.02e-11
+ mcm4d_ca_w_0_300_s_3_300 = 1.07e-05  mcm4d_cc_w_0_300_s_3_300 = 2.65e-11  mcm4d_cf_w_0_300_s_3_300 = 1.44e-11
+ mcm4d_ca_w_0_300_s_9_000 = 1.07e-05  mcm4d_cc_w_0_300_s_9_000 = 8.78e-12  mcm4d_cf_w_0_300_s_9_000 = 2.66e-11
+ mcm4d_ca_w_2_400_s_0_300 = 1.07e-05  mcm4d_cc_w_2_400_s_0_300 = 1.50e-10  mcm4d_cf_w_2_400_s_0_300 = 1.44e-12
+ mcm4d_ca_w_2_400_s_0_360 = 1.07e-05  mcm4d_cc_w_2_400_s_0_360 = 1.40e-10  mcm4d_cf_w_2_400_s_0_360 = 1.76e-12
+ mcm4d_ca_w_2_400_s_0_450 = 1.07e-05  mcm4d_cc_w_2_400_s_0_450 = 1.27e-10  mcm4d_cf_w_2_400_s_0_450 = 2.23e-12
+ mcm4d_ca_w_2_400_s_0_600 = 1.07e-05  mcm4d_cc_w_2_400_s_0_600 = 1.09e-10  mcm4d_cf_w_2_400_s_0_600 = 3.00e-12
+ mcm4d_ca_w_2_400_s_0_800 = 1.07e-05  mcm4d_cc_w_2_400_s_0_800 = 9.31e-11  mcm4d_cf_w_2_400_s_0_800 = 4.00e-12
+ mcm4d_ca_w_2_400_s_1_000 = 1.07e-05  mcm4d_cc_w_2_400_s_1_000 = 8.10e-11  mcm4d_cf_w_2_400_s_1_000 = 4.99e-12
+ mcm4d_ca_w_2_400_s_1_200 = 1.07e-05  mcm4d_cc_w_2_400_s_1_200 = 7.19e-11  mcm4d_cf_w_2_400_s_1_200 = 5.96e-12
+ mcm4d_ca_w_2_400_s_2_100 = 1.07e-05  mcm4d_cc_w_2_400_s_2_100 = 4.94e-11  mcm4d_cf_w_2_400_s_2_100 = 1.00e-11
+ mcm4d_ca_w_2_400_s_3_300 = 1.07e-05  mcm4d_cc_w_2_400_s_3_300 = 3.53e-11  mcm4d_cf_w_2_400_s_3_300 = 1.48e-11
+ mcm4d_ca_w_2_400_s_9_000 = 1.07e-05  mcm4d_cc_w_2_400_s_9_000 = 1.29e-11  mcm4d_cf_w_2_400_s_9_000 = 2.88e-11
+ mcm4p1_ca_w_0_300_s_0_300 = 1.17e-05  mcm4p1_cc_w_0_300_s_0_300 = 1.21e-10  mcm4p1_cf_w_0_300_s_0_300 = 1.55e-12
+ mcm4p1_ca_w_0_300_s_0_360 = 1.17e-05  mcm4p1_cc_w_0_300_s_0_360 = 1.12e-10  mcm4p1_cf_w_0_300_s_0_360 = 1.90e-12
+ mcm4p1_ca_w_0_300_s_0_450 = 1.17e-05  mcm4p1_cc_w_0_300_s_0_450 = 1.00e-10  mcm4p1_cf_w_0_300_s_0_450 = 2.43e-12
+ mcm4p1_ca_w_0_300_s_0_600 = 1.17e-05  mcm4p1_cc_w_0_300_s_0_600 = 8.61e-11  mcm4p1_cf_w_0_300_s_0_600 = 3.29e-12
+ mcm4p1_ca_w_0_300_s_0_800 = 1.17e-05  mcm4p1_cc_w_0_300_s_0_800 = 7.27e-11  mcm4p1_cf_w_0_300_s_0_800 = 4.33e-12
+ mcm4p1_ca_w_0_300_s_1_000 = 1.17e-05  mcm4p1_cc_w_0_300_s_1_000 = 6.26e-11  mcm4p1_cf_w_0_300_s_1_000 = 5.39e-12
+ mcm4p1_ca_w_0_300_s_1_200 = 1.17e-05  mcm4p1_cc_w_0_300_s_1_200 = 5.52e-11  mcm4p1_cf_w_0_300_s_1_200 = 6.43e-12
+ mcm4p1_ca_w_0_300_s_2_100 = 1.17e-05  mcm4p1_cc_w_0_300_s_2_100 = 3.67e-11  mcm4p1_cf_w_0_300_s_2_100 = 1.10e-11
+ mcm4p1_ca_w_0_300_s_3_300 = 1.17e-05  mcm4p1_cc_w_0_300_s_3_300 = 2.58e-11  mcm4p1_cf_w_0_300_s_3_300 = 1.55e-11
+ mcm4p1_ca_w_0_300_s_9_000 = 1.17e-05  mcm4p1_cc_w_0_300_s_9_000 = 8.23e-12  mcm4p1_cf_w_0_300_s_9_000 = 2.79e-11
+ mcm4p1_ca_w_2_400_s_0_300 = 1.17e-05  mcm4p1_cc_w_2_400_s_0_300 = 1.49e-10  mcm4p1_cf_w_2_400_s_0_300 = 1.59e-12
+ mcm4p1_ca_w_2_400_s_0_360 = 1.17e-05  mcm4p1_cc_w_2_400_s_0_360 = 1.39e-10  mcm4p1_cf_w_2_400_s_0_360 = 1.94e-12
+ mcm4p1_ca_w_2_400_s_0_450 = 1.17e-05  mcm4p1_cc_w_2_400_s_0_450 = 1.26e-10  mcm4p1_cf_w_2_400_s_0_450 = 2.45e-12
+ mcm4p1_ca_w_2_400_s_0_600 = 1.17e-05  mcm4p1_cc_w_2_400_s_0_600 = 1.09e-10  mcm4p1_cf_w_2_400_s_0_600 = 3.29e-12
+ mcm4p1_ca_w_2_400_s_0_800 = 1.17e-05  mcm4p1_cc_w_2_400_s_0_800 = 9.22e-11  mcm4p1_cf_w_2_400_s_0_800 = 4.39e-12
+ mcm4p1_ca_w_2_400_s_1_000 = 1.17e-05  mcm4p1_cc_w_2_400_s_1_000 = 8.01e-11  mcm4p1_cf_w_2_400_s_1_000 = 5.47e-12
+ mcm4p1_ca_w_2_400_s_1_200 = 1.17e-05  mcm4p1_cc_w_2_400_s_1_200 = 7.10e-11  mcm4p1_cf_w_2_400_s_1_200 = 6.52e-12
+ mcm4p1_ca_w_2_400_s_2_100 = 1.17e-05  mcm4p1_cc_w_2_400_s_2_100 = 4.85e-11  mcm4p1_cf_w_2_400_s_2_100 = 1.09e-11
+ mcm4p1_ca_w_2_400_s_3_300 = 1.17e-05  mcm4p1_cc_w_2_400_s_3_300 = 3.44e-11  mcm4p1_cf_w_2_400_s_3_300 = 1.60e-11
+ mcm4p1_ca_w_2_400_s_9_000 = 1.17e-05  mcm4p1_cc_w_2_400_s_9_000 = 1.22e-11  mcm4p1_cf_w_2_400_s_9_000 = 3.04e-11
+ mcm4l1_ca_w_0_300_s_0_300 = 1.34e-05  mcm4l1_cc_w_0_300_s_0_300 = 1.20e-10  mcm4l1_cf_w_0_300_s_0_300 = 1.76e-12
+ mcm4l1_ca_w_0_300_s_0_360 = 1.34e-05  mcm4l1_cc_w_0_300_s_0_360 = 1.11e-10  mcm4l1_cf_w_0_300_s_0_360 = 2.14e-12
+ mcm4l1_ca_w_0_300_s_0_450 = 1.34e-05  mcm4l1_cc_w_0_300_s_0_450 = 9.97e-11  mcm4l1_cf_w_0_300_s_0_450 = 2.74e-12
+ mcm4l1_ca_w_0_300_s_0_600 = 1.34e-05  mcm4l1_cc_w_0_300_s_0_600 = 8.56e-11  mcm4l1_cf_w_0_300_s_0_600 = 3.72e-12
+ mcm4l1_ca_w_0_300_s_0_800 = 1.34e-05  mcm4l1_cc_w_0_300_s_0_800 = 7.20e-11  mcm4l1_cf_w_0_300_s_0_800 = 4.89e-12
+ mcm4l1_ca_w_0_300_s_1_000 = 1.34e-05  mcm4l1_cc_w_0_300_s_1_000 = 6.18e-11  mcm4l1_cf_w_0_300_s_1_000 = 6.07e-12
+ mcm4l1_ca_w_0_300_s_1_200 = 1.34e-05  mcm4l1_cc_w_0_300_s_1_200 = 5.43e-11  mcm4l1_cf_w_0_300_s_1_200 = 7.23e-12
+ mcm4l1_ca_w_0_300_s_2_100 = 1.34e-05  mcm4l1_cc_w_0_300_s_2_100 = 3.57e-11  mcm4l1_cf_w_0_300_s_2_100 = 1.23e-11
+ mcm4l1_ca_w_0_300_s_3_300 = 1.34e-05  mcm4l1_cc_w_0_300_s_3_300 = 2.47e-11  mcm4l1_cf_w_0_300_s_3_300 = 1.72e-11
+ mcm4l1_ca_w_0_300_s_9_000 = 1.34e-05  mcm4l1_cc_w_0_300_s_9_000 = 7.47e-12  mcm4l1_cf_w_0_300_s_9_000 = 2.98e-11
+ mcm4l1_ca_w_2_400_s_0_300 = 1.34e-05  mcm4l1_cc_w_2_400_s_0_300 = 1.48e-10  mcm4l1_cf_w_2_400_s_0_300 = 1.77e-12
+ mcm4l1_ca_w_2_400_s_0_360 = 1.34e-05  mcm4l1_cc_w_2_400_s_0_360 = 1.38e-10  mcm4l1_cf_w_2_400_s_0_360 = 2.16e-12
+ mcm4l1_ca_w_2_400_s_0_450 = 1.34e-05  mcm4l1_cc_w_2_400_s_0_450 = 1.25e-10  mcm4l1_cf_w_2_400_s_0_450 = 2.74e-12
+ mcm4l1_ca_w_2_400_s_0_600 = 1.34e-05  mcm4l1_cc_w_2_400_s_0_600 = 1.07e-10  mcm4l1_cf_w_2_400_s_0_600 = 3.69e-12
+ mcm4l1_ca_w_2_400_s_0_800 = 1.34e-05  mcm4l1_cc_w_2_400_s_0_800 = 9.10e-11  mcm4l1_cf_w_2_400_s_0_800 = 4.93e-12
+ mcm4l1_ca_w_2_400_s_1_000 = 1.34e-05  mcm4l1_cc_w_2_400_s_1_000 = 7.88e-11  mcm4l1_cf_w_2_400_s_1_000 = 6.14e-12
+ mcm4l1_ca_w_2_400_s_1_200 = 1.34e-05  mcm4l1_cc_w_2_400_s_1_200 = 6.98e-11  mcm4l1_cf_w_2_400_s_1_200 = 7.30e-12
+ mcm4l1_ca_w_2_400_s_2_100 = 1.34e-05  mcm4l1_cc_w_2_400_s_2_100 = 4.72e-11  mcm4l1_cf_w_2_400_s_2_100 = 1.21e-11
+ mcm4l1_ca_w_2_400_s_3_300 = 1.34e-05  mcm4l1_cc_w_2_400_s_3_300 = 3.31e-11  mcm4l1_cf_w_2_400_s_3_300 = 1.76e-11
+ mcm4l1_ca_w_2_400_s_9_000 = 1.34e-05  mcm4l1_cc_w_2_400_s_9_000 = 1.13e-11  mcm4l1_cf_w_2_400_s_9_000 = 3.25e-11
+ mcm4m1_ca_w_0_300_s_0_300 = 1.73e-05  mcm4m1_cc_w_0_300_s_0_300 = 1.19e-10  mcm4m1_cf_w_0_300_s_0_300 = 2.27e-12
+ mcm4m1_ca_w_0_300_s_0_360 = 1.73e-05  mcm4m1_cc_w_0_300_s_0_360 = 1.10e-10  mcm4m1_cf_w_0_300_s_0_360 = 2.76e-12
+ mcm4m1_ca_w_0_300_s_0_450 = 1.73e-05  mcm4m1_cc_w_0_300_s_0_450 = 9.86e-11  mcm4m1_cf_w_0_300_s_0_450 = 3.52e-12
+ mcm4m1_ca_w_0_300_s_0_600 = 1.73e-05  mcm4m1_cc_w_0_300_s_0_600 = 8.43e-11  mcm4m1_cf_w_0_300_s_0_600 = 4.75e-12
+ mcm4m1_ca_w_0_300_s_0_800 = 1.73e-05  mcm4m1_cc_w_0_300_s_0_800 = 7.04e-11  mcm4m1_cf_w_0_300_s_0_800 = 6.24e-12
+ mcm4m1_ca_w_0_300_s_1_000 = 1.73e-05  mcm4m1_cc_w_0_300_s_1_000 = 6.02e-11  mcm4m1_cf_w_0_300_s_1_000 = 7.74e-12
+ mcm4m1_ca_w_0_300_s_1_200 = 1.73e-05  mcm4m1_cc_w_0_300_s_1_200 = 5.25e-11  mcm4m1_cf_w_0_300_s_1_200 = 9.17e-12
+ mcm4m1_ca_w_0_300_s_2_100 = 1.73e-05  mcm4m1_cc_w_0_300_s_2_100 = 3.35e-11  mcm4m1_cf_w_0_300_s_2_100 = 1.52e-11
+ mcm4m1_ca_w_0_300_s_3_300 = 1.73e-05  mcm4m1_cc_w_0_300_s_3_300 = 2.25e-11  mcm4m1_cf_w_0_300_s_3_300 = 2.09e-11
+ mcm4m1_ca_w_0_300_s_9_000 = 1.73e-05  mcm4m1_cc_w_0_300_s_9_000 = 6.17e-12  mcm4m1_cf_w_0_300_s_9_000 = 3.37e-11
+ mcm4m1_ca_w_2_400_s_0_300 = 1.73e-05  mcm4m1_cc_w_2_400_s_0_300 = 1.45e-10  mcm4m1_cf_w_2_400_s_0_300 = 2.27e-12
+ mcm4m1_ca_w_2_400_s_0_360 = 1.73e-05  mcm4m1_cc_w_2_400_s_0_360 = 1.35e-10  mcm4m1_cf_w_2_400_s_0_360 = 2.77e-12
+ mcm4m1_ca_w_2_400_s_0_450 = 1.73e-05  mcm4m1_cc_w_2_400_s_0_450 = 1.22e-10  mcm4m1_cf_w_2_400_s_0_450 = 3.51e-12
+ mcm4m1_ca_w_2_400_s_0_600 = 1.73e-05  mcm4m1_cc_w_2_400_s_0_600 = 1.04e-10  mcm4m1_cf_w_2_400_s_0_600 = 4.71e-12
+ mcm4m1_ca_w_2_400_s_0_800 = 1.73e-05  mcm4m1_cc_w_2_400_s_0_800 = 8.84e-11  mcm4m1_cf_w_2_400_s_0_800 = 6.27e-12
+ mcm4m1_ca_w_2_400_s_1_000 = 1.73e-05  mcm4m1_cc_w_2_400_s_1_000 = 7.61e-11  mcm4m1_cf_w_2_400_s_1_000 = 7.80e-12
+ mcm4m1_ca_w_2_400_s_1_200 = 1.73e-05  mcm4m1_cc_w_2_400_s_1_200 = 6.71e-11  mcm4m1_cf_w_2_400_s_1_200 = 9.24e-12
+ mcm4m1_ca_w_2_400_s_2_100 = 1.73e-05  mcm4m1_cc_w_2_400_s_2_100 = 4.46e-11  mcm4m1_cf_w_2_400_s_2_100 = 1.51e-11
+ mcm4m1_ca_w_2_400_s_3_300 = 1.73e-05  mcm4m1_cc_w_2_400_s_3_300 = 3.06e-11  mcm4m1_cf_w_2_400_s_3_300 = 2.15e-11
+ mcm4m1_ca_w_2_400_s_9_000 = 1.73e-05  mcm4m1_cc_w_2_400_s_9_000 = 9.75e-12  mcm4m1_cf_w_2_400_s_9_000 = 3.68e-11
+ mcm4m2_ca_w_0_300_s_0_300 = 2.38e-05  mcm4m2_cc_w_0_300_s_0_300 = 1.18e-10  mcm4m2_cf_w_0_300_s_0_300 = 3.09e-12
+ mcm4m2_ca_w_0_300_s_0_360 = 2.38e-05  mcm4m2_cc_w_0_300_s_0_360 = 1.09e-10  mcm4m2_cf_w_0_300_s_0_360 = 3.76e-12
+ mcm4m2_ca_w_0_300_s_0_450 = 2.38e-05  mcm4m2_cc_w_0_300_s_0_450 = 9.72e-11  mcm4m2_cf_w_0_300_s_0_450 = 4.76e-12
+ mcm4m2_ca_w_0_300_s_0_600 = 2.38e-05  mcm4m2_cc_w_0_300_s_0_600 = 8.22e-11  mcm4m2_cf_w_0_300_s_0_600 = 6.39e-12
+ mcm4m2_ca_w_0_300_s_0_800 = 2.38e-05  mcm4m2_cc_w_0_300_s_0_800 = 6.82e-11  mcm4m2_cf_w_0_300_s_0_800 = 8.38e-12
+ mcm4m2_ca_w_0_300_s_1_000 = 2.38e-05  mcm4m2_cc_w_0_300_s_1_000 = 5.79e-11  mcm4m2_cf_w_0_300_s_1_000 = 1.03e-11
+ mcm4m2_ca_w_0_300_s_1_200 = 2.38e-05  mcm4m2_cc_w_0_300_s_1_200 = 5.01e-11  mcm4m2_cf_w_0_300_s_1_200 = 1.22e-11
+ mcm4m2_ca_w_0_300_s_2_100 = 2.38e-05  mcm4m2_cc_w_0_300_s_2_100 = 3.07e-11  mcm4m2_cf_w_0_300_s_2_100 = 1.96e-11
+ mcm4m2_ca_w_0_300_s_3_300 = 2.38e-05  mcm4m2_cc_w_0_300_s_3_300 = 1.98e-11  mcm4m2_cf_w_0_300_s_3_300 = 2.60e-11
+ mcm4m2_ca_w_0_300_s_9_000 = 2.38e-05  mcm4m2_cc_w_0_300_s_9_000 = 4.88e-12  mcm4m2_cf_w_0_300_s_9_000 = 3.85e-11
+ mcm4m2_ca_w_2_400_s_0_300 = 2.38e-05  mcm4m2_cc_w_2_400_s_0_300 = 1.42e-10  mcm4m2_cf_w_2_400_s_0_300 = 3.09e-12
+ mcm4m2_ca_w_2_400_s_0_360 = 2.38e-05  mcm4m2_cc_w_2_400_s_0_360 = 1.32e-10  mcm4m2_cf_w_2_400_s_0_360 = 3.76e-12
+ mcm4m2_ca_w_2_400_s_0_450 = 2.38e-05  mcm4m2_cc_w_2_400_s_0_450 = 1.18e-10  mcm4m2_cf_w_2_400_s_0_450 = 4.75e-12
+ mcm4m2_ca_w_2_400_s_0_600 = 2.38e-05  mcm4m2_cc_w_2_400_s_0_600 = 1.01e-10  mcm4m2_cf_w_2_400_s_0_600 = 6.36e-12
+ mcm4m2_ca_w_2_400_s_0_800 = 2.38e-05  mcm4m2_cc_w_2_400_s_0_800 = 8.50e-11  mcm4m2_cf_w_2_400_s_0_800 = 8.42e-12
+ mcm4m2_ca_w_2_400_s_1_000 = 2.38e-05  mcm4m2_cc_w_2_400_s_1_000 = 7.27e-11  mcm4m2_cf_w_2_400_s_1_000 = 1.04e-11
+ mcm4m2_ca_w_2_400_s_1_200 = 2.38e-05  mcm4m2_cc_w_2_400_s_1_200 = 6.36e-11  mcm4m2_cf_w_2_400_s_1_200 = 1.22e-11
+ mcm4m2_ca_w_2_400_s_2_100 = 2.38e-05  mcm4m2_cc_w_2_400_s_2_100 = 4.14e-11  mcm4m2_cf_w_2_400_s_2_100 = 1.95e-11
+ mcm4m2_ca_w_2_400_s_3_300 = 2.38e-05  mcm4m2_cc_w_2_400_s_3_300 = 2.77e-11  mcm4m2_cf_w_2_400_s_3_300 = 2.68e-11
+ mcm4m2_ca_w_2_400_s_9_000 = 2.38e-05  mcm4m2_cc_w_2_400_s_9_000 = 8.20e-12  mcm4m2_cf_w_2_400_s_9_000 = 4.23e-11
+ mcm4m3_ca_w_0_300_s_0_300 = 1.42e-04  mcm4m3_cc_w_0_300_s_0_300 = 1.02e-10  mcm4m3_cf_w_0_300_s_0_300 = 1.61e-11
+ mcm4m3_ca_w_0_300_s_0_360 = 1.42e-04  mcm4m3_cc_w_0_300_s_0_360 = 9.28e-11  mcm4m3_cf_w_0_300_s_0_360 = 1.90e-11
+ mcm4m3_ca_w_0_300_s_0_450 = 1.42e-04  mcm4m3_cc_w_0_300_s_0_450 = 8.12e-11  mcm4m3_cf_w_0_300_s_0_450 = 2.29e-11
+ mcm4m3_ca_w_0_300_s_0_600 = 1.42e-04  mcm4m3_cc_w_0_300_s_0_600 = 6.63e-11  mcm4m3_cf_w_0_300_s_0_600 = 2.86e-11
+ mcm4m3_ca_w_0_300_s_0_800 = 1.42e-04  mcm4m3_cc_w_0_300_s_0_800 = 5.27e-11  mcm4m3_cf_w_0_300_s_0_800 = 3.44e-11
+ mcm4m3_ca_w_0_300_s_1_000 = 1.42e-04  mcm4m3_cc_w_0_300_s_1_000 = 4.28e-11  mcm4m3_cf_w_0_300_s_1_000 = 3.92e-11
+ mcm4m3_ca_w_0_300_s_1_200 = 1.42e-04  mcm4m3_cc_w_0_300_s_1_200 = 3.56e-11  mcm4m3_cf_w_0_300_s_1_200 = 4.31e-11
+ mcm4m3_ca_w_0_300_s_2_100 = 1.42e-04  mcm4m3_cc_w_0_300_s_2_100 = 1.84e-11  mcm4m3_cf_w_0_300_s_2_100 = 5.51e-11
+ mcm4m3_ca_w_0_300_s_3_300 = 1.42e-04  mcm4m3_cc_w_0_300_s_3_300 = 1.05e-11  mcm4m3_cf_w_0_300_s_3_300 = 6.18e-11
+ mcm4m3_ca_w_0_300_s_9_000 = 1.42e-04  mcm4m3_cc_w_0_300_s_9_000 = 2.05e-12  mcm4m3_cf_w_0_300_s_9_000 = 7.01e-11
+ mcm4m3_ca_w_2_400_s_0_300 = 1.42e-04  mcm4m3_cc_w_2_400_s_0_300 = 1.23e-10  mcm4m3_cf_w_2_400_s_0_300 = 1.60e-11
+ mcm4m3_ca_w_2_400_s_0_360 = 1.42e-04  mcm4m3_cc_w_2_400_s_0_360 = 1.13e-10  mcm4m3_cf_w_2_400_s_0_360 = 1.90e-11
+ mcm4m3_ca_w_2_400_s_0_450 = 1.42e-04  mcm4m3_cc_w_2_400_s_0_450 = 9.98e-11  mcm4m3_cf_w_2_400_s_0_450 = 2.29e-11
+ mcm4m3_ca_w_2_400_s_0_600 = 1.42e-04  mcm4m3_cc_w_2_400_s_0_600 = 8.34e-11  mcm4m3_cf_w_2_400_s_0_600 = 2.85e-11
+ mcm4m3_ca_w_2_400_s_0_800 = 1.42e-04  mcm4m3_cc_w_2_400_s_0_800 = 6.78e-11  mcm4m3_cf_w_2_400_s_0_800 = 3.44e-11
+ mcm4m3_ca_w_2_400_s_1_000 = 1.42e-04  mcm4m3_cc_w_2_400_s_1_000 = 5.67e-11  mcm4m3_cf_w_2_400_s_1_000 = 3.93e-11
+ mcm4m3_ca_w_2_400_s_1_200 = 1.42e-04  mcm4m3_cc_w_2_400_s_1_200 = 4.85e-11  mcm4m3_cf_w_2_400_s_1_200 = 4.32e-11
+ mcm4m3_ca_w_2_400_s_2_100 = 1.42e-04  mcm4m3_cc_w_2_400_s_2_100 = 2.91e-11  mcm4m3_cf_w_2_400_s_2_100 = 5.52e-11
+ mcm4m3_ca_w_2_400_s_3_300 = 1.42e-04  mcm4m3_cc_w_2_400_s_3_300 = 1.79e-11  mcm4m3_cf_w_2_400_s_3_300 = 6.41e-11
+ mcm4m3_ca_w_2_400_s_9_000 = 1.42e-04  mcm4m3_cc_w_2_400_s_9_000 = 4.40e-12  mcm4m3_cf_w_2_400_s_9_000 = 7.68e-11
+ mcm5f_ca_w_1_600_s_1_600 = 7.33e-06  mcm5f_cc_w_1_600_s_1_600 = 8.49e-11  mcm5f_cf_w_1_600_s_1_600 = 5.39e-12
+ mcm5f_ca_w_1_600_s_1_700 = 7.33e-06  mcm5f_cc_w_1_600_s_1_700 = 8.06e-11  mcm5f_cf_w_1_600_s_1_700 = 5.73e-12
+ mcm5f_ca_w_1_600_s_1_900 = 7.33e-06  mcm5f_cc_w_1_600_s_1_900 = 7.29e-11  mcm5f_cf_w_1_600_s_1_900 = 6.40e-12
+ mcm5f_ca_w_1_600_s_2_000 = 7.33e-06  mcm5f_cc_w_1_600_s_2_000 = 6.98e-11  mcm5f_cf_w_1_600_s_2_000 = 6.72e-12
+ mcm5f_ca_w_1_600_s_2_400 = 7.33e-06  mcm5f_cc_w_1_600_s_2_400 = 5.98e-11  mcm5f_cf_w_1_600_s_2_400 = 8.02e-12
+ mcm5f_ca_w_1_600_s_2_800 = 7.33e-06  mcm5f_cc_w_1_600_s_2_800 = 5.26e-11  mcm5f_cf_w_1_600_s_2_800 = 9.30e-12
+ mcm5f_ca_w_1_600_s_3_200 = 7.33e-06  mcm5f_cc_w_1_600_s_3_200 = 4.70e-11  mcm5f_cf_w_1_600_s_3_200 = 1.05e-11
+ mcm5f_ca_w_1_600_s_4_800 = 7.33e-06  mcm5f_cc_w_1_600_s_4_800 = 3.31e-11  mcm5f_cf_w_1_600_s_4_800 = 1.50e-11
+ mcm5f_ca_w_1_600_s_10_000 = 7.33e-06  mcm5f_cc_w_1_600_s_10_000 = 1.54e-11  mcm5f_cf_w_1_600_s_10_000 = 2.53e-11
+ mcm5f_ca_w_1_600_s_12_000 = 7.33e-06  mcm5f_cc_w_1_600_s_12_000 = 1.22e-11  mcm5f_cf_w_1_600_s_12_000 = 2.78e-11
+ mcm5f_ca_w_4_000_s_1_600 = 7.33e-06  mcm5f_cc_w_4_000_s_1_600 = 9.22e-11  mcm5f_cf_w_4_000_s_1_600 = 5.39e-12
+ mcm5f_ca_w_4_000_s_1_700 = 7.33e-06  mcm5f_cc_w_4_000_s_1_700 = 8.75e-11  mcm5f_cf_w_4_000_s_1_700 = 5.73e-12
+ mcm5f_ca_w_4_000_s_1_900 = 7.33e-06  mcm5f_cc_w_4_000_s_1_900 = 7.97e-11  mcm5f_cf_w_4_000_s_1_900 = 6.40e-12
+ mcm5f_ca_w_4_000_s_2_000 = 7.33e-06  mcm5f_cc_w_4_000_s_2_000 = 7.64e-11  mcm5f_cf_w_4_000_s_2_000 = 6.73e-12
+ mcm5f_ca_w_4_000_s_2_400 = 7.33e-06  mcm5f_cc_w_4_000_s_2_400 = 6.58e-11  mcm5f_cf_w_4_000_s_2_400 = 8.04e-12
+ mcm5f_ca_w_4_000_s_2_800 = 7.33e-06  mcm5f_cc_w_4_000_s_2_800 = 5.80e-11  mcm5f_cf_w_4_000_s_2_800 = 9.31e-12
+ mcm5f_ca_w_4_000_s_3_200 = 7.33e-06  mcm5f_cc_w_4_000_s_3_200 = 5.21e-11  mcm5f_cf_w_4_000_s_3_200 = 1.05e-11
+ mcm5f_ca_w_4_000_s_4_800 = 7.33e-06  mcm5f_cc_w_4_000_s_4_800 = 3.72e-11  mcm5f_cf_w_4_000_s_4_800 = 1.51e-11
+ mcm5f_ca_w_4_000_s_10_000 = 7.33e-06  mcm5f_cc_w_4_000_s_10_000 = 1.81e-11  mcm5f_cf_w_4_000_s_10_000 = 2.57e-11
+ mcm5f_ca_w_4_000_s_12_000 = 7.33e-06  mcm5f_cc_w_4_000_s_12_000 = 1.46e-11  mcm5f_cf_w_4_000_s_12_000 = 2.84e-11
+ mcm5d_ca_w_1_600_s_1_600 = 7.72e-06  mcm5d_cc_w_1_600_s_1_600 = 8.45e-11  mcm5d_cf_w_1_600_s_1_600 = 5.67e-12
+ mcm5d_ca_w_1_600_s_1_700 = 7.72e-06  mcm5d_cc_w_1_600_s_1_700 = 8.03e-11  mcm5d_cf_w_1_600_s_1_700 = 6.02e-12
+ mcm5d_ca_w_1_600_s_1_900 = 7.72e-06  mcm5d_cc_w_1_600_s_1_900 = 7.25e-11  mcm5d_cf_w_1_600_s_1_900 = 6.72e-12
+ mcm5d_ca_w_1_600_s_2_000 = 7.72e-06  mcm5d_cc_w_1_600_s_2_000 = 6.94e-11  mcm5d_cf_w_1_600_s_2_000 = 7.07e-12
+ mcm5d_ca_w_1_600_s_2_400 = 7.72e-06  mcm5d_cc_w_1_600_s_2_400 = 5.94e-11  mcm5d_cf_w_1_600_s_2_400 = 8.43e-12
+ mcm5d_ca_w_1_600_s_2_800 = 7.72e-06  mcm5d_cc_w_1_600_s_2_800 = 5.21e-11  mcm5d_cf_w_1_600_s_2_800 = 9.76e-12
+ mcm5d_ca_w_1_600_s_3_200 = 7.72e-06  mcm5d_cc_w_1_600_s_3_200 = 4.65e-11  mcm5d_cf_w_1_600_s_3_200 = 1.10e-11
+ mcm5d_ca_w_1_600_s_4_800 = 7.72e-06  mcm5d_cc_w_1_600_s_4_800 = 3.26e-11  mcm5d_cf_w_1_600_s_4_800 = 1.57e-11
+ mcm5d_ca_w_1_600_s_10_000 = 7.72e-06  mcm5d_cc_w_1_600_s_10_000 = 1.49e-11  mcm5d_cf_w_1_600_s_10_000 = 2.62e-11
+ mcm5d_ca_w_1_600_s_12_000 = 7.72e-06  mcm5d_cc_w_1_600_s_12_000 = 1.18e-11  mcm5d_cf_w_1_600_s_12_000 = 2.87e-11
+ mcm5d_ca_w_4_000_s_1_600 = 7.72e-06  mcm5d_cc_w_4_000_s_1_600 = 9.17e-11  mcm5d_cf_w_4_000_s_1_600 = 5.67e-12
+ mcm5d_ca_w_4_000_s_1_700 = 7.72e-06  mcm5d_cc_w_4_000_s_1_700 = 8.70e-11  mcm5d_cf_w_4_000_s_1_700 = 6.03e-12
+ mcm5d_ca_w_4_000_s_1_900 = 7.72e-06  mcm5d_cc_w_4_000_s_1_900 = 7.91e-11  mcm5d_cf_w_4_000_s_1_900 = 6.73e-12
+ mcm5d_ca_w_4_000_s_2_000 = 7.72e-06  mcm5d_cc_w_4_000_s_2_000 = 7.58e-11  mcm5d_cf_w_4_000_s_2_000 = 7.08e-12
+ mcm5d_ca_w_4_000_s_2_400 = 7.72e-06  mcm5d_cc_w_4_000_s_2_400 = 6.52e-11  mcm5d_cf_w_4_000_s_2_400 = 8.44e-12
+ mcm5d_ca_w_4_000_s_2_800 = 7.72e-06  mcm5d_cc_w_4_000_s_2_800 = 5.75e-11  mcm5d_cf_w_4_000_s_2_800 = 9.78e-12
+ mcm5d_ca_w_4_000_s_3_200 = 7.72e-06  mcm5d_cc_w_4_000_s_3_200 = 5.16e-11  mcm5d_cf_w_4_000_s_3_200 = 1.11e-11
+ mcm5d_ca_w_4_000_s_4_800 = 7.72e-06  mcm5d_cc_w_4_000_s_4_800 = 3.67e-11  mcm5d_cf_w_4_000_s_4_800 = 1.58e-11
+ mcm5d_ca_w_4_000_s_10_000 = 7.72e-06  mcm5d_cc_w_4_000_s_10_000 = 1.76e-11  mcm5d_cf_w_4_000_s_10_000 = 2.66e-11
+ mcm5d_ca_w_4_000_s_12_000 = 7.72e-06  mcm5d_cc_w_4_000_s_12_000 = 1.42e-11  mcm5d_cf_w_4_000_s_12_000 = 2.94e-11
+ mcm5p1_ca_w_1_600_s_1_600 = 8.24e-06  mcm5p1_cc_w_1_600_s_1_600 = 8.41e-11  mcm5p1_cf_w_1_600_s_1_600 = 6.03e-12
+ mcm5p1_ca_w_1_600_s_1_700 = 8.24e-06  mcm5p1_cc_w_1_600_s_1_700 = 7.97e-11  mcm5p1_cf_w_1_600_s_1_700 = 6.41e-12
+ mcm5p1_ca_w_1_600_s_1_900 = 8.24e-06  mcm5p1_cc_w_1_600_s_1_900 = 7.19e-11  mcm5p1_cf_w_1_600_s_1_900 = 7.15e-12
+ mcm5p1_ca_w_1_600_s_2_000 = 8.24e-06  mcm5p1_cc_w_1_600_s_2_000 = 6.89e-11  mcm5p1_cf_w_1_600_s_2_000 = 7.52e-12
+ mcm5p1_ca_w_1_600_s_2_400 = 8.24e-06  mcm5p1_cc_w_1_600_s_2_400 = 5.88e-11  mcm5p1_cf_w_1_600_s_2_400 = 8.96e-12
+ mcm5p1_ca_w_1_600_s_2_800 = 8.24e-06  mcm5p1_cc_w_1_600_s_2_800 = 5.15e-11  mcm5p1_cf_w_1_600_s_2_800 = 1.04e-11
+ mcm5p1_ca_w_1_600_s_3_200 = 8.24e-06  mcm5p1_cc_w_1_600_s_3_200 = 4.59e-11  mcm5p1_cf_w_1_600_s_3_200 = 1.17e-11
+ mcm5p1_ca_w_1_600_s_4_800 = 8.24e-06  mcm5p1_cc_w_1_600_s_4_800 = 3.20e-11  mcm5p1_cf_w_1_600_s_4_800 = 1.66e-11
+ mcm5p1_ca_w_1_600_s_10_000 = 8.24e-06  mcm5p1_cc_w_1_600_s_10_000 = 1.44e-11  mcm5p1_cf_w_1_600_s_10_000 = 2.73e-11
+ mcm5p1_ca_w_1_600_s_12_000 = 8.24e-06  mcm5p1_cc_w_1_600_s_12_000 = 1.13e-11  mcm5p1_cf_w_1_600_s_12_000 = 2.99e-11
+ mcm5p1_ca_w_4_000_s_1_600 = 8.24e-06  mcm5p1_cc_w_4_000_s_1_600 = 9.10e-11  mcm5p1_cf_w_4_000_s_1_600 = 6.05e-12
+ mcm5p1_ca_w_4_000_s_1_700 = 8.24e-06  mcm5p1_cc_w_4_000_s_1_700 = 8.63e-11  mcm5p1_cf_w_4_000_s_1_700 = 6.42e-12
+ mcm5p1_ca_w_4_000_s_1_900 = 8.24e-06  mcm5p1_cc_w_4_000_s_1_900 = 7.84e-11  mcm5p1_cf_w_4_000_s_1_900 = 7.16e-12
+ mcm5p1_ca_w_4_000_s_2_000 = 8.24e-06  mcm5p1_cc_w_4_000_s_2_000 = 7.51e-11  mcm5p1_cf_w_4_000_s_2_000 = 7.53e-12
+ mcm5p1_ca_w_4_000_s_2_400 = 8.24e-06  mcm5p1_cc_w_4_000_s_2_400 = 6.45e-11  mcm5p1_cf_w_4_000_s_2_400 = 8.98e-12
+ mcm5p1_ca_w_4_000_s_2_800 = 8.24e-06  mcm5p1_cc_w_4_000_s_2_800 = 5.68e-11  mcm5p1_cf_w_4_000_s_2_800 = 1.04e-11
+ mcm5p1_ca_w_4_000_s_3_200 = 8.24e-06  mcm5p1_cc_w_4_000_s_3_200 = 5.09e-11  mcm5p1_cf_w_4_000_s_3_200 = 1.17e-11
+ mcm5p1_ca_w_4_000_s_4_800 = 8.24e-06  mcm5p1_cc_w_4_000_s_4_800 = 3.60e-11  mcm5p1_cf_w_4_000_s_4_800 = 1.66e-11
+ mcm5p1_ca_w_4_000_s_10_000 = 8.24e-06  mcm5p1_cc_w_4_000_s_10_000 = 1.71e-11  mcm5p1_cf_w_4_000_s_10_000 = 2.78e-11
+ mcm5p1_ca_w_4_000_s_12_000 = 8.24e-06  mcm5p1_cc_w_4_000_s_12_000 = 1.37e-11  mcm5p1_cf_w_4_000_s_12_000 = 3.05e-11
+ mcm5l1_ca_w_1_600_s_1_600 = 8.99e-06  mcm5l1_cc_w_1_600_s_1_600 = 8.35e-11  mcm5l1_cf_w_1_600_s_1_600 = 6.55e-12
+ mcm5l1_ca_w_1_600_s_1_700 = 8.99e-06  mcm5l1_cc_w_1_600_s_1_700 = 7.90e-11  mcm5l1_cf_w_1_600_s_1_700 = 6.96e-12
+ mcm5l1_ca_w_1_600_s_1_900 = 8.99e-06  mcm5l1_cc_w_1_600_s_1_900 = 7.12e-11  mcm5l1_cf_w_1_600_s_1_900 = 7.76e-12
+ mcm5l1_ca_w_1_600_s_2_000 = 8.99e-06  mcm5l1_cc_w_1_600_s_2_000 = 6.82e-11  mcm5l1_cf_w_1_600_s_2_000 = 8.16e-12
+ mcm5l1_ca_w_1_600_s_2_400 = 8.99e-06  mcm5l1_cc_w_1_600_s_2_400 = 5.80e-11  mcm5l1_cf_w_1_600_s_2_400 = 9.71e-12
+ mcm5l1_ca_w_1_600_s_2_800 = 8.99e-06  mcm5l1_cc_w_1_600_s_2_800 = 5.07e-11  mcm5l1_cf_w_1_600_s_2_800 = 1.12e-11
+ mcm5l1_ca_w_1_600_s_3_200 = 8.99e-06  mcm5l1_cc_w_1_600_s_3_200 = 4.51e-11  mcm5l1_cf_w_1_600_s_3_200 = 1.26e-11
+ mcm5l1_ca_w_1_600_s_4_800 = 8.99e-06  mcm5l1_cc_w_1_600_s_4_800 = 3.11e-11  mcm5l1_cf_w_1_600_s_4_800 = 1.78e-11
+ mcm5l1_ca_w_1_600_s_10_000 = 8.99e-06  mcm5l1_cc_w_1_600_s_10_000 = 1.37e-11  mcm5l1_cf_w_1_600_s_10_000 = 2.89e-11
+ mcm5l1_ca_w_1_600_s_12_000 = 8.99e-06  mcm5l1_cc_w_1_600_s_12_000 = 1.06e-11  mcm5l1_cf_w_1_600_s_12_000 = 3.14e-11
+ mcm5l1_ca_w_4_000_s_1_600 = 8.99e-06  mcm5l1_cc_w_4_000_s_1_600 = 9.04e-11  mcm5l1_cf_w_4_000_s_1_600 = 6.56e-12
+ mcm5l1_ca_w_4_000_s_1_700 = 8.99e-06  mcm5l1_cc_w_4_000_s_1_700 = 8.55e-11  mcm5l1_cf_w_4_000_s_1_700 = 6.96e-12
+ mcm5l1_ca_w_4_000_s_1_900 = 8.99e-06  mcm5l1_cc_w_4_000_s_1_900 = 7.75e-11  mcm5l1_cf_w_4_000_s_1_900 = 7.77e-12
+ mcm5l1_ca_w_4_000_s_2_000 = 8.99e-06  mcm5l1_cc_w_4_000_s_2_000 = 7.42e-11  mcm5l1_cf_w_4_000_s_2_000 = 8.16e-12
+ mcm5l1_ca_w_4_000_s_2_400 = 8.99e-06  mcm5l1_cc_w_4_000_s_2_400 = 6.36e-11  mcm5l1_cf_w_4_000_s_2_400 = 9.73e-12
+ mcm5l1_ca_w_4_000_s_2_800 = 8.99e-06  mcm5l1_cc_w_4_000_s_2_800 = 5.59e-11  mcm5l1_cf_w_4_000_s_2_800 = 1.12e-11
+ mcm5l1_ca_w_4_000_s_3_200 = 8.99e-06  mcm5l1_cc_w_4_000_s_3_200 = 4.99e-11  mcm5l1_cf_w_4_000_s_3_200 = 1.27e-11
+ mcm5l1_ca_w_4_000_s_4_800 = 8.99e-06  mcm5l1_cc_w_4_000_s_4_800 = 3.51e-11  mcm5l1_cf_w_4_000_s_4_800 = 1.79e-11
+ mcm5l1_ca_w_4_000_s_10_000 = 8.99e-06  mcm5l1_cc_w_4_000_s_10_000 = 1.63e-11  mcm5l1_cf_w_4_000_s_10_000 = 2.94e-11
+ mcm5l1_ca_w_4_000_s_12_000 = 8.99e-06  mcm5l1_cc_w_4_000_s_12_000 = 1.30e-11  mcm5l1_cf_w_4_000_s_12_000 = 3.21e-11
+ mcm5m1_ca_w_1_600_s_1_600 = 1.06e-05  mcm5m1_cc_w_1_600_s_1_600 = 8.20e-11  mcm5m1_cf_w_1_600_s_1_600 = 7.68e-12
+ mcm5m1_ca_w_1_600_s_1_700 = 1.06e-05  mcm5m1_cc_w_1_600_s_1_700 = 7.74e-11  mcm5m1_cf_w_1_600_s_1_700 = 8.15e-12
+ mcm5m1_ca_w_1_600_s_1_900 = 1.06e-05  mcm5m1_cc_w_1_600_s_1_900 = 6.97e-11  mcm5m1_cf_w_1_600_s_1_900 = 9.08e-12
+ mcm5m1_ca_w_1_600_s_2_000 = 1.06e-05  mcm5m1_cc_w_1_600_s_2_000 = 6.66e-11  mcm5m1_cf_w_1_600_s_2_000 = 9.53e-12
+ mcm5m1_ca_w_1_600_s_2_400 = 1.06e-05  mcm5m1_cc_w_1_600_s_2_400 = 5.64e-11  mcm5m1_cf_w_1_600_s_2_400 = 1.13e-11
+ mcm5m1_ca_w_1_600_s_2_800 = 1.06e-05  mcm5m1_cc_w_1_600_s_2_800 = 4.91e-11  mcm5m1_cf_w_1_600_s_2_800 = 1.30e-11
+ mcm5m1_ca_w_1_600_s_3_200 = 1.06e-05  mcm5m1_cc_w_1_600_s_3_200 = 4.35e-11  mcm5m1_cf_w_1_600_s_3_200 = 1.47e-11
+ mcm5m1_ca_w_1_600_s_4_800 = 1.06e-05  mcm5m1_cc_w_1_600_s_4_800 = 2.95e-11  mcm5m1_cf_w_1_600_s_4_800 = 2.04e-11
+ mcm5m1_ca_w_1_600_s_10_000 = 1.06e-05  mcm5m1_cc_w_1_600_s_10_000 = 1.24e-11  mcm5m1_cf_w_1_600_s_10_000 = 3.20e-11
+ mcm5m1_ca_w_1_600_s_12_000 = 1.06e-05  mcm5m1_cc_w_1_600_s_12_000 = 9.53e-12  mcm5m1_cf_w_1_600_s_12_000 = 3.45e-11
+ mcm5m1_ca_w_4_000_s_1_600 = 1.06e-05  mcm5m1_cc_w_4_000_s_1_600 = 8.86e-11  mcm5m1_cf_w_4_000_s_1_600 = 7.67e-12
+ mcm5m1_ca_w_4_000_s_1_700 = 1.06e-05  mcm5m1_cc_w_4_000_s_1_700 = 8.37e-11  mcm5m1_cf_w_4_000_s_1_700 = 8.15e-12
+ mcm5m1_ca_w_4_000_s_1_900 = 1.06e-05  mcm5m1_cc_w_4_000_s_1_900 = 7.58e-11  mcm5m1_cf_w_4_000_s_1_900 = 9.08e-12
+ mcm5m1_ca_w_4_000_s_2_000 = 1.06e-05  mcm5m1_cc_w_4_000_s_2_000 = 7.25e-11  mcm5m1_cf_w_4_000_s_2_000 = 9.54e-12
+ mcm5m1_ca_w_4_000_s_2_400 = 1.06e-05  mcm5m1_cc_w_4_000_s_2_400 = 6.18e-11  mcm5m1_cf_w_4_000_s_2_400 = 1.13e-11
+ mcm5m1_ca_w_4_000_s_2_800 = 1.06e-05  mcm5m1_cc_w_4_000_s_2_800 = 5.41e-11  mcm5m1_cf_w_4_000_s_2_800 = 1.30e-11
+ mcm5m1_ca_w_4_000_s_3_200 = 1.06e-05  mcm5m1_cc_w_4_000_s_3_200 = 4.82e-11  mcm5m1_cf_w_4_000_s_3_200 = 1.47e-11
+ mcm5m1_ca_w_4_000_s_4_800 = 1.06e-05  mcm5m1_cc_w_4_000_s_4_800 = 3.34e-11  mcm5m1_cf_w_4_000_s_4_800 = 2.05e-11
+ mcm5m1_ca_w_4_000_s_10_000 = 1.06e-05  mcm5m1_cc_w_4_000_s_10_000 = 1.50e-11  mcm5m1_cf_w_4_000_s_10_000 = 3.26e-11
+ mcm5m1_ca_w_4_000_s_12_000 = 1.06e-05  mcm5m1_cc_w_4_000_s_12_000 = 1.18e-11  mcm5m1_cf_w_4_000_s_12_000 = 3.53e-11
+ mcm5m2_ca_w_1_600_s_1_600 = 1.27e-05  mcm5m2_cc_w_1_600_s_1_600 = 8.03e-11  mcm5m2_cf_w_1_600_s_1_600 = 9.11e-12
+ mcm5m2_ca_w_1_600_s_1_700 = 1.27e-05  mcm5m2_cc_w_1_600_s_1_700 = 7.57e-11  mcm5m2_cf_w_1_600_s_1_700 = 9.66e-12
+ mcm5m2_ca_w_1_600_s_1_900 = 1.27e-05  mcm5m2_cc_w_1_600_s_1_900 = 6.81e-11  mcm5m2_cf_w_1_600_s_1_900 = 1.07e-11
+ mcm5m2_ca_w_1_600_s_2_000 = 1.27e-05  mcm5m2_cc_w_1_600_s_2_000 = 6.49e-11  mcm5m2_cf_w_1_600_s_2_000 = 1.13e-11
+ mcm5m2_ca_w_1_600_s_2_400 = 1.27e-05  mcm5m2_cc_w_1_600_s_2_400 = 5.47e-11  mcm5m2_cf_w_1_600_s_2_400 = 1.33e-11
+ mcm5m2_ca_w_1_600_s_2_800 = 1.27e-05  mcm5m2_cc_w_1_600_s_2_800 = 4.73e-11  mcm5m2_cf_w_1_600_s_2_800 = 1.53e-11
+ mcm5m2_ca_w_1_600_s_3_200 = 1.27e-05  mcm5m2_cc_w_1_600_s_3_200 = 4.17e-11  mcm5m2_cf_w_1_600_s_3_200 = 1.72e-11
+ mcm5m2_ca_w_1_600_s_4_800 = 1.27e-05  mcm5m2_cc_w_1_600_s_4_800 = 2.77e-11  mcm5m2_cf_w_1_600_s_4_800 = 2.36e-11
+ mcm5m2_ca_w_1_600_s_10_000 = 1.27e-05  mcm5m2_cc_w_1_600_s_10_000 = 1.11e-11  mcm5m2_cf_w_1_600_s_10_000 = 3.56e-11
+ mcm5m2_ca_w_1_600_s_12_000 = 1.27e-05  mcm5m2_cc_w_1_600_s_12_000 = 8.40e-12  mcm5m2_cf_w_1_600_s_12_000 = 3.79e-11
+ mcm5m2_ca_w_4_000_s_1_600 = 1.27e-05  mcm5m2_cc_w_4_000_s_1_600 = 8.67e-11  mcm5m2_cf_w_4_000_s_1_600 = 9.10e-12
+ mcm5m2_ca_w_4_000_s_1_700 = 1.27e-05  mcm5m2_cc_w_4_000_s_1_700 = 8.18e-11  mcm5m2_cf_w_4_000_s_1_700 = 9.65e-12
+ mcm5m2_ca_w_4_000_s_1_900 = 1.27e-05  mcm5m2_cc_w_4_000_s_1_900 = 7.39e-11  mcm5m2_cf_w_4_000_s_1_900 = 1.07e-11
+ mcm5m2_ca_w_4_000_s_2_000 = 1.27e-05  mcm5m2_cc_w_4_000_s_2_000 = 7.06e-11  mcm5m2_cf_w_4_000_s_2_000 = 1.13e-11
+ mcm5m2_ca_w_4_000_s_2_400 = 1.27e-05  mcm5m2_cc_w_4_000_s_2_400 = 5.99e-11  mcm5m2_cf_w_4_000_s_2_400 = 1.33e-11
+ mcm5m2_ca_w_4_000_s_2_800 = 1.27e-05  mcm5m2_cc_w_4_000_s_2_800 = 5.22e-11  mcm5m2_cf_w_4_000_s_2_800 = 1.53e-11
+ mcm5m2_ca_w_4_000_s_3_200 = 1.27e-05  mcm5m2_cc_w_4_000_s_3_200 = 4.63e-11  mcm5m2_cf_w_4_000_s_3_200 = 1.72e-11
+ mcm5m2_ca_w_4_000_s_4_800 = 1.27e-05  mcm5m2_cc_w_4_000_s_4_800 = 3.16e-11  mcm5m2_cf_w_4_000_s_4_800 = 2.37e-11
+ mcm5m2_ca_w_4_000_s_10_000 = 1.27e-05  mcm5m2_cc_w_4_000_s_10_000 = 1.36e-11  mcm5m2_cf_w_4_000_s_10_000 = 3.62e-11
+ mcm5m2_ca_w_4_000_s_12_000 = 1.27e-05  mcm5m2_cc_w_4_000_s_12_000 = 1.06e-11  mcm5m2_cf_w_4_000_s_12_000 = 3.88e-11
+ mcm5m3_ca_w_1_600_s_1_600 = 2.30e-05  mcm5m3_cc_w_1_600_s_1_600 = 7.40e-11  mcm5m3_cf_w_1_600_s_1_600 = 1.56e-11
+ mcm5m3_ca_w_1_600_s_1_700 = 2.30e-05  mcm5m3_cc_w_1_600_s_1_700 = 6.95e-11  mcm5m3_cf_w_1_600_s_1_700 = 1.65e-11
+ mcm5m3_ca_w_1_600_s_1_900 = 2.30e-05  mcm5m3_cc_w_1_600_s_1_900 = 6.18e-11  mcm5m3_cf_w_1_600_s_1_900 = 1.82e-11
+ mcm5m3_ca_w_1_600_s_2_000 = 2.30e-05  mcm5m3_cc_w_1_600_s_2_000 = 5.87e-11  mcm5m3_cf_w_1_600_s_2_000 = 1.90e-11
+ mcm5m3_ca_w_1_600_s_2_400 = 2.30e-05  mcm5m3_cc_w_1_600_s_2_400 = 4.86e-11  mcm5m3_cf_w_1_600_s_2_400 = 2.22e-11
+ mcm5m3_ca_w_1_600_s_2_800 = 2.30e-05  mcm5m3_cc_w_1_600_s_2_800 = 4.12e-11  mcm5m3_cf_w_1_600_s_2_800 = 2.51e-11
+ mcm5m3_ca_w_1_600_s_3_200 = 2.30e-05  mcm5m3_cc_w_1_600_s_3_200 = 3.57e-11  mcm5m3_cf_w_1_600_s_3_200 = 2.76e-11
+ mcm5m3_ca_w_1_600_s_4_800 = 2.30e-05  mcm5m3_cc_w_1_600_s_4_800 = 2.22e-11  mcm5m3_cf_w_1_600_s_4_800 = 3.58e-11
+ mcm5m3_ca_w_1_600_s_10_000 = 2.30e-05  mcm5m3_cc_w_1_600_s_10_000 = 7.80e-12  mcm5m3_cf_w_1_600_s_10_000 = 4.78e-11
+ mcm5m3_ca_w_1_600_s_12_000 = 2.30e-05  mcm5m3_cc_w_1_600_s_12_000 = 5.80e-12  mcm5m3_cf_w_1_600_s_12_000 = 4.97e-11
+ mcm5m3_ca_w_4_000_s_1_600 = 2.30e-05  mcm5m3_cc_w_4_000_s_1_600 = 7.99e-11  mcm5m3_cf_w_4_000_s_1_600 = 1.56e-11
+ mcm5m3_ca_w_4_000_s_1_700 = 2.30e-05  mcm5m3_cc_w_4_000_s_1_700 = 7.51e-11  mcm5m3_cf_w_4_000_s_1_700 = 1.65e-11
+ mcm5m3_ca_w_4_000_s_1_900 = 2.30e-05  mcm5m3_cc_w_4_000_s_1_900 = 6.75e-11  mcm5m3_cf_w_4_000_s_1_900 = 1.82e-11
+ mcm5m3_ca_w_4_000_s_2_000 = 2.30e-05  mcm5m3_cc_w_4_000_s_2_000 = 6.41e-11  mcm5m3_cf_w_4_000_s_2_000 = 1.90e-11
+ mcm5m3_ca_w_4_000_s_2_400 = 2.30e-05  mcm5m3_cc_w_4_000_s_2_400 = 5.35e-11  mcm5m3_cf_w_4_000_s_2_400 = 2.22e-11
+ mcm5m3_ca_w_4_000_s_2_800 = 2.30e-05  mcm5m3_cc_w_4_000_s_2_800 = 4.60e-11  mcm5m3_cf_w_4_000_s_2_800 = 2.51e-11
+ mcm5m3_ca_w_4_000_s_3_200 = 2.30e-05  mcm5m3_cc_w_4_000_s_3_200 = 4.02e-11  mcm5m3_cf_w_4_000_s_3_200 = 2.77e-11
+ mcm5m3_ca_w_4_000_s_4_800 = 2.30e-05  mcm5m3_cc_w_4_000_s_4_800 = 2.61e-11  mcm5m3_cf_w_4_000_s_4_800 = 3.60e-11
+ mcm5m3_ca_w_4_000_s_10_000 = 2.30e-05  mcm5m3_cc_w_4_000_s_10_000 = 1.03e-11  mcm5m3_cf_w_4_000_s_10_000 = 4.88e-11
+ mcm5m3_ca_w_4_000_s_12_000 = 2.30e-05  mcm5m3_cc_w_4_000_s_12_000 = 7.85e-12  mcm5m3_cf_w_4_000_s_12_000 = 5.10e-11
+ mcm5m4_ca_w_1_600_s_1_600 = 9.63e-05  mcm5m4_cc_w_1_600_s_1_600 = 5.93e-11  mcm5m4_cf_w_1_600_s_1_600 = 4.69e-11
+ mcm5m4_ca_w_1_600_s_1_700 = 9.63e-05  mcm5m4_cc_w_1_600_s_1_700 = 5.48e-11  mcm5m4_cf_w_1_600_s_1_700 = 4.87e-11
+ mcm5m4_ca_w_1_600_s_1_900 = 9.63e-05  mcm5m4_cc_w_1_600_s_1_900 = 4.75e-11  mcm5m4_cf_w_1_600_s_1_900 = 5.21e-11
+ mcm5m4_ca_w_1_600_s_2_000 = 9.63e-05  mcm5m4_cc_w_1_600_s_2_000 = 4.45e-11  mcm5m4_cf_w_1_600_s_2_000 = 5.36e-11
+ mcm5m4_ca_w_1_600_s_2_400 = 9.63e-05  mcm5m4_cc_w_1_600_s_2_400 = 3.53e-11  mcm5m4_cf_w_1_600_s_2_400 = 5.88e-11
+ mcm5m4_ca_w_1_600_s_2_800 = 9.63e-05  mcm5m4_cc_w_1_600_s_2_800 = 2.89e-11  mcm5m4_cf_w_1_600_s_2_800 = 6.31e-11
+ mcm5m4_ca_w_1_600_s_3_200 = 9.63e-05  mcm5m4_cc_w_1_600_s_3_200 = 2.42e-11  mcm5m4_cf_w_1_600_s_3_200 = 6.64e-11
+ mcm5m4_ca_w_1_600_s_4_800 = 9.63e-05  mcm5m4_cc_w_1_600_s_4_800 = 1.37e-11  mcm5m4_cf_w_1_600_s_4_800 = 7.50e-11
+ mcm5m4_ca_w_1_600_s_10_000 = 9.63e-05  mcm5m4_cc_w_1_600_s_10_000 = 4.35e-12  mcm5m4_cf_w_1_600_s_10_000 = 8.40e-11
+ mcm5m4_ca_w_1_600_s_12_000 = 9.63e-05  mcm5m4_cc_w_1_600_s_12_000 = 3.25e-12  mcm5m4_cf_w_1_600_s_12_000 = 8.52e-11
+ mcm5m4_ca_w_4_000_s_1_600 = 9.63e-05  mcm5m4_cc_w_4_000_s_1_600 = 6.52e-11  mcm5m4_cf_w_4_000_s_1_600 = 4.69e-11
+ mcm5m4_ca_w_4_000_s_1_700 = 9.63e-05  mcm5m4_cc_w_4_000_s_1_700 = 6.06e-11  mcm5m4_cf_w_4_000_s_1_700 = 4.87e-11
+ mcm5m4_ca_w_4_000_s_1_900 = 9.63e-05  mcm5m4_cc_w_4_000_s_1_900 = 5.31e-11  mcm5m4_cf_w_4_000_s_1_900 = 5.21e-11
+ mcm5m4_ca_w_4_000_s_2_000 = 9.63e-05  mcm5m4_cc_w_4_000_s_2_000 = 5.00e-11  mcm5m4_cf_w_4_000_s_2_000 = 5.36e-11
+ mcm5m4_ca_w_4_000_s_2_400 = 9.63e-05  mcm5m4_cc_w_4_000_s_2_400 = 4.03e-11  mcm5m4_cf_w_4_000_s_2_400 = 5.88e-11
+ mcm5m4_ca_w_4_000_s_2_800 = 9.63e-05  mcm5m4_cc_w_4_000_s_2_800 = 3.38e-11  mcm5m4_cf_w_4_000_s_2_800 = 6.31e-11
+ mcm5m4_ca_w_4_000_s_3_200 = 9.63e-05  mcm5m4_cc_w_4_000_s_3_200 = 2.89e-11  mcm5m4_cf_w_4_000_s_3_200 = 6.66e-11
+ mcm5m4_ca_w_4_000_s_4_800 = 9.63e-05  mcm5m4_cc_w_4_000_s_4_800 = 1.76e-11  mcm5m4_cf_w_4_000_s_4_800 = 7.55e-11
+ mcm5m4_ca_w_4_000_s_10_000 = 9.63e-05  mcm5m4_cc_w_4_000_s_10_000 = 6.55e-12  mcm5m4_cf_w_4_000_s_10_000 = 8.59e-11
+ mcm5m4_ca_w_4_000_s_12_000 = 9.63e-05  mcm5m4_cc_w_4_000_s_12_000 = 5.00e-12  mcm5m4_cf_w_4_000_s_12_000 = 8.74e-11
+ mcrdlf_ca_w_10_000_s_5_000 = 3.26e-06  mcrdlf_cc_w_10_000_s_5_000 = 6.41e-11  mcrdlf_cf_w_10_000_s_5_000 = 6.52e-12
+ mcrdlf_ca_w_10_000_s_8_000 = 3.26e-06  mcrdlf_cc_w_10_000_s_8_000 = 4.43e-11  mcrdlf_cf_w_10_000_s_8_000 = 1.04e-11
+ mcrdlf_ca_w_10_000_s_10_000 = 3.26e-06  mcrdlf_cc_w_10_000_s_10_000 = 3.71e-11  mcrdlf_cf_w_10_000_s_10_000 = 1.27e-11
+ mcrdlf_ca_w_10_000_s_12_000 = 3.26e-06  mcrdlf_cc_w_10_000_s_12_000 = 3.21e-11  mcrdlf_cf_w_10_000_s_12_000 = 1.48e-11
+ mcrdlf_ca_w_10_000_s_30_000 = 3.26e-06  mcrdlf_cc_w_10_000_s_30_000 = 1.33e-11  mcrdlf_cf_w_10_000_s_30_000 = 2.68e-11
+ mcrdlf_ca_w_40_000_s_5_000 = 3.26e-06  mcrdlf_cc_w_40_000_s_5_000 = 7.56e-11  mcrdlf_cf_w_40_000_s_5_000 = 6.60e-12
+ mcrdlf_ca_w_40_000_s_8_000 = 3.26e-06  mcrdlf_cc_w_40_000_s_8_000 = 5.48e-11  mcrdlf_cf_w_40_000_s_8_000 = 1.05e-11
+ mcrdlf_ca_w_40_000_s_10_000 = 3.26e-06  mcrdlf_cc_w_40_000_s_10_000 = 4.71e-11  mcrdlf_cf_w_40_000_s_10_000 = 1.28e-11
+ mcrdlf_ca_w_40_000_s_12_000 = 3.26e-06  mcrdlf_cc_w_40_000_s_12_000 = 4.15e-11  mcrdlf_cf_w_40_000_s_12_000 = 1.49e-11
+ mcrdlf_ca_w_40_000_s_30_000 = 3.26e-06  mcrdlf_cc_w_40_000_s_30_000 = 2.05e-11  mcrdlf_cf_w_40_000_s_30_000 = 2.75e-11
+ mcrdld_ca_w_10_000_s_5_000 = 3.34e-06  mcrdld_cc_w_10_000_s_5_000 = 6.39e-11  mcrdld_cf_w_10_000_s_5_000 = 6.66e-12
+ mcrdld_ca_w_10_000_s_8_000 = 3.34e-06  mcrdld_cc_w_10_000_s_8_000 = 4.41e-11  mcrdld_cf_w_10_000_s_8_000 = 1.06e-11
+ mcrdld_ca_w_10_000_s_10_000 = 3.34e-06  mcrdld_cc_w_10_000_s_10_000 = 3.69e-11  mcrdld_cf_w_10_000_s_10_000 = 1.29e-11
+ mcrdld_ca_w_10_000_s_12_000 = 3.34e-06  mcrdld_cc_w_10_000_s_12_000 = 3.18e-11  mcrdld_cf_w_10_000_s_12_000 = 1.51e-11
+ mcrdld_ca_w_10_000_s_30_000 = 3.34e-06  mcrdld_cc_w_10_000_s_30_000 = 1.31e-11  mcrdld_cf_w_10_000_s_30_000 = 2.72e-11
+ mcrdld_ca_w_40_000_s_5_000 = 3.34e-06  mcrdld_cc_w_40_000_s_5_000 = 7.54e-11  mcrdld_cf_w_40_000_s_5_000 = 6.75e-12
+ mcrdld_ca_w_40_000_s_8_000 = 3.34e-06  mcrdld_cc_w_40_000_s_8_000 = 5.45e-11  mcrdld_cf_w_40_000_s_8_000 = 1.07e-11
+ mcrdld_ca_w_40_000_s_10_000 = 3.34e-06  mcrdld_cc_w_40_000_s_10_000 = 4.68e-11  mcrdld_cf_w_40_000_s_10_000 = 1.30e-11
+ mcrdld_ca_w_40_000_s_12_000 = 3.34e-06  mcrdld_cc_w_40_000_s_12_000 = 4.13e-11  mcrdld_cf_w_40_000_s_12_000 = 1.52e-11
+ mcrdld_ca_w_40_000_s_30_000 = 3.34e-06  mcrdld_cc_w_40_000_s_30_000 = 2.03e-11  mcrdld_cf_w_40_000_s_30_000 = 2.78e-11
+ mcrdlp1_ca_w_10_000_s_5_000 = 3.43e-06  mcrdlp1_cc_w_10_000_s_5_000 = 6.36e-11  mcrdlp1_cf_w_10_000_s_5_000 = 6.83e-12
+ mcrdlp1_ca_w_10_000_s_8_000 = 3.43e-06  mcrdlp1_cc_w_10_000_s_8_000 = 4.38e-11  mcrdlp1_cf_w_10_000_s_8_000 = 1.09e-11
+ mcrdlp1_ca_w_10_000_s_10_000 = 3.43e-06  mcrdlp1_cc_w_10_000_s_10_000 = 3.67e-11  mcrdlp1_cf_w_10_000_s_10_000 = 1.32e-11
+ mcrdlp1_ca_w_10_000_s_12_000 = 3.43e-06  mcrdlp1_cc_w_10_000_s_12_000 = 3.16e-11  mcrdlp1_cf_w_10_000_s_12_000 = 1.54e-11
+ mcrdlp1_ca_w_10_000_s_30_000 = 3.43e-06  mcrdlp1_cc_w_10_000_s_30_000 = 1.30e-11  mcrdlp1_cf_w_10_000_s_30_000 = 2.76e-11
+ mcrdlp1_ca_w_40_000_s_5_000 = 3.43e-06  mcrdlp1_cc_w_40_000_s_5_000 = 7.51e-11  mcrdlp1_cf_w_40_000_s_5_000 = 6.91e-12
+ mcrdlp1_ca_w_40_000_s_8_000 = 3.43e-06  mcrdlp1_cc_w_40_000_s_8_000 = 5.42e-11  mcrdlp1_cf_w_40_000_s_8_000 = 1.09e-11
+ mcrdlp1_ca_w_40_000_s_10_000 = 3.43e-06  mcrdlp1_cc_w_40_000_s_10_000 = 4.65e-11  mcrdlp1_cf_w_40_000_s_10_000 = 1.33e-11
+ mcrdlp1_ca_w_40_000_s_12_000 = 3.43e-06  mcrdlp1_cc_w_40_000_s_12_000 = 4.10e-11  mcrdlp1_cf_w_40_000_s_12_000 = 1.55e-11
+ mcrdlp1_ca_w_40_000_s_30_000 = 3.43e-06  mcrdlp1_cc_w_40_000_s_30_000 = 2.01e-11  mcrdlp1_cf_w_40_000_s_30_000 = 2.82e-11
+ mcrdll1_ca_w_10_000_s_5_000 = 3.55e-06  mcrdll1_cc_w_10_000_s_5_000 = 6.33e-11  mcrdll1_cf_w_10_000_s_5_000 = 7.05e-12
+ mcrdll1_ca_w_10_000_s_8_000 = 3.55e-06  mcrdll1_cc_w_10_000_s_8_000 = 4.35e-11  mcrdll1_cf_w_10_000_s_8_000 = 1.12e-11
+ mcrdll1_ca_w_10_000_s_10_000 = 3.55e-06  mcrdll1_cc_w_10_000_s_10_000 = 3.63e-11  mcrdll1_cf_w_10_000_s_10_000 = 1.36e-11
+ mcrdll1_ca_w_10_000_s_12_000 = 3.55e-06  mcrdll1_cc_w_10_000_s_12_000 = 3.12e-11  mcrdll1_cf_w_10_000_s_12_000 = 1.58e-11
+ mcrdll1_ca_w_10_000_s_30_000 = 3.55e-06  mcrdll1_cc_w_10_000_s_30_000 = 1.27e-11  mcrdll1_cf_w_10_000_s_30_000 = 2.80e-11
+ mcrdll1_ca_w_40_000_s_5_000 = 3.55e-06  mcrdll1_cc_w_40_000_s_5_000 = 7.48e-11  mcrdll1_cf_w_40_000_s_5_000 = 7.12e-12
+ mcrdll1_ca_w_40_000_s_8_000 = 3.55e-06  mcrdll1_cc_w_40_000_s_8_000 = 5.39e-11  mcrdll1_cf_w_40_000_s_8_000 = 1.12e-11
+ mcrdll1_ca_w_40_000_s_10_000 = 3.55e-06  mcrdll1_cc_w_40_000_s_10_000 = 4.62e-11  mcrdll1_cf_w_40_000_s_10_000 = 1.37e-11
+ mcrdll1_ca_w_40_000_s_12_000 = 3.55e-06  mcrdll1_cc_w_40_000_s_12_000 = 4.06e-11  mcrdll1_cf_w_40_000_s_12_000 = 1.59e-11
+ mcrdll1_ca_w_40_000_s_30_000 = 3.55e-06  mcrdll1_cc_w_40_000_s_30_000 = 1.99e-11  mcrdll1_cf_w_40_000_s_30_000 = 2.88e-11
+ mcrdlm1_ca_w_10_000_s_5_000 = 3.79e-06  mcrdlm1_cc_w_10_000_s_5_000 = 6.27e-11  mcrdlm1_cf_w_10_000_s_5_000 = 7.45e-12
+ mcrdlm1_ca_w_10_000_s_8_000 = 3.79e-06  mcrdlm1_cc_w_10_000_s_8_000 = 4.28e-11  mcrdlm1_cf_w_10_000_s_8_000 = 1.18e-11
+ mcrdlm1_ca_w_10_000_s_10_000 = 3.79e-06  mcrdlm1_cc_w_10_000_s_10_000 = 3.57e-11  mcrdlm1_cf_w_10_000_s_10_000 = 1.43e-11
+ mcrdlm1_ca_w_10_000_s_12_000 = 3.79e-06  mcrdlm1_cc_w_10_000_s_12_000 = 3.07e-11  mcrdlm1_cf_w_10_000_s_12_000 = 1.66e-11
+ mcrdlm1_ca_w_10_000_s_30_000 = 3.79e-06  mcrdlm1_cc_w_10_000_s_30_000 = 1.24e-11  mcrdlm1_cf_w_10_000_s_30_000 = 2.89e-11
+ mcrdlm1_ca_w_40_000_s_5_000 = 3.79e-06  mcrdlm1_cc_w_40_000_s_5_000 = 7.41e-11  mcrdlm1_cf_w_40_000_s_5_000 = 7.51e-12
+ mcrdlm1_ca_w_40_000_s_8_000 = 3.79e-06  mcrdlm1_cc_w_40_000_s_8_000 = 5.33e-11  mcrdlm1_cf_w_40_000_s_8_000 = 1.18e-11
+ mcrdlm1_ca_w_40_000_s_10_000 = 3.79e-06  mcrdlm1_cc_w_40_000_s_10_000 = 4.56e-11  mcrdlm1_cf_w_40_000_s_10_000 = 1.44e-11
+ mcrdlm1_ca_w_40_000_s_12_000 = 3.79e-06  mcrdlm1_cc_w_40_000_s_12_000 = 4.01e-11  mcrdlm1_cf_w_40_000_s_12_000 = 1.66e-11
+ mcrdlm1_ca_w_40_000_s_30_000 = 3.79e-06  mcrdlm1_cc_w_40_000_s_30_000 = 1.94e-11  mcrdlm1_cf_w_40_000_s_30_000 = 2.97e-11
+ mcrdlm2_ca_w_10_000_s_5_000 = 4.02e-06  mcrdlm2_cc_w_10_000_s_5_000 = 6.20e-11  mcrdlm2_cf_w_10_000_s_5_000 = 7.88e-12
+ mcrdlm2_ca_w_10_000_s_8_000 = 4.02e-06  mcrdlm2_cc_w_10_000_s_8_000 = 4.23e-11  mcrdlm2_cf_w_10_000_s_8_000 = 1.24e-11
+ mcrdlm2_ca_w_10_000_s_10_000 = 4.02e-06  mcrdlm2_cc_w_10_000_s_10_000 = 3.51e-11  mcrdlm2_cf_w_10_000_s_10_000 = 1.50e-11
+ mcrdlm2_ca_w_10_000_s_12_000 = 4.02e-06  mcrdlm2_cc_w_10_000_s_12_000 = 3.01e-11  mcrdlm2_cf_w_10_000_s_12_000 = 1.73e-11
+ mcrdlm2_ca_w_10_000_s_30_000 = 4.02e-06  mcrdlm2_cc_w_10_000_s_30_000 = 1.21e-11  mcrdlm2_cf_w_10_000_s_30_000 = 2.98e-11
+ mcrdlm2_ca_w_40_000_s_5_000 = 4.02e-06  mcrdlm2_cc_w_40_000_s_5_000 = 7.35e-11  mcrdlm2_cf_w_40_000_s_5_000 = 7.94e-12
+ mcrdlm2_ca_w_40_000_s_8_000 = 4.02e-06  mcrdlm2_cc_w_40_000_s_8_000 = 5.27e-11  mcrdlm2_cf_w_40_000_s_8_000 = 1.24e-11
+ mcrdlm2_ca_w_40_000_s_10_000 = 4.02e-06  mcrdlm2_cc_w_40_000_s_10_000 = 4.51e-11  mcrdlm2_cf_w_40_000_s_10_000 = 1.51e-11
+ mcrdlm2_ca_w_40_000_s_12_000 = 4.02e-06  mcrdlm2_cc_w_40_000_s_12_000 = 3.96e-11  mcrdlm2_cf_w_40_000_s_12_000 = 1.74e-11
+ mcrdlm2_ca_w_40_000_s_30_000 = 4.02e-06  mcrdlm2_cc_w_40_000_s_30_000 = 1.91e-11  mcrdlm2_cf_w_40_000_s_30_000 = 3.06e-11
+ mcrdlm3_ca_w_10_000_s_5_000 = 4.69e-06  mcrdlm3_cc_w_10_000_s_5_000 = 6.05e-11  mcrdlm3_cf_w_10_000_s_5_000 = 8.99e-12
+ mcrdlm3_ca_w_10_000_s_8_000 = 4.69e-06  mcrdlm3_cc_w_10_000_s_8_000 = 4.08e-11  mcrdlm3_cf_w_10_000_s_8_000 = 1.40e-11
+ mcrdlm3_ca_w_10_000_s_10_000 = 4.69e-06  mcrdlm3_cc_w_10_000_s_10_000 = 3.38e-11  mcrdlm3_cf_w_10_000_s_10_000 = 1.68e-11
+ mcrdlm3_ca_w_10_000_s_12_000 = 4.69e-06  mcrdlm3_cc_w_10_000_s_12_000 = 2.88e-11  mcrdlm3_cf_w_10_000_s_12_000 = 1.93e-11
+ mcrdlm3_ca_w_10_000_s_30_000 = 4.69e-06  mcrdlm3_cc_w_10_000_s_30_000 = 1.12e-11  mcrdlm3_cf_w_10_000_s_30_000 = 3.19e-11
+ mcrdlm3_ca_w_40_000_s_5_000 = 4.69e-06  mcrdlm3_cc_w_40_000_s_5_000 = 7.20e-11  mcrdlm3_cf_w_40_000_s_5_000 = 8.98e-12
+ mcrdlm3_ca_w_40_000_s_8_000 = 4.69e-06  mcrdlm3_cc_w_40_000_s_8_000 = 5.13e-11  mcrdlm3_cf_w_40_000_s_8_000 = 1.40e-11
+ mcrdlm3_ca_w_40_000_s_10_000 = 4.69e-06  mcrdlm3_cc_w_40_000_s_10_000 = 4.37e-11  mcrdlm3_cf_w_40_000_s_10_000 = 1.68e-11
+ mcrdlm3_ca_w_40_000_s_12_000 = 4.69e-06  mcrdlm3_cc_w_40_000_s_12_000 = 3.83e-11  mcrdlm3_cf_w_40_000_s_12_000 = 1.93e-11
+ mcrdlm3_ca_w_40_000_s_30_000 = 4.69e-06  mcrdlm3_cc_w_40_000_s_30_000 = 1.83e-11  mcrdlm3_cf_w_40_000_s_30_000 = 3.28e-11
+ mcrdlm4_ca_w_10_000_s_5_000 = 5.55e-06  mcrdlm4_cc_w_10_000_s_5_000 = 5.89e-11  mcrdlm4_cf_w_10_000_s_5_000 = 1.04e-11
+ mcrdlm4_ca_w_10_000_s_8_000 = 5.55e-06  mcrdlm4_cc_w_10_000_s_8_000 = 3.93e-11  mcrdlm4_cf_w_10_000_s_8_000 = 1.59e-11
+ mcrdlm4_ca_w_10_000_s_10_000 = 5.55e-06  mcrdlm4_cc_w_10_000_s_10_000 = 3.23e-11  mcrdlm4_cf_w_10_000_s_10_000 = 1.89e-11
+ mcrdlm4_ca_w_10_000_s_12_000 = 5.55e-06  mcrdlm4_cc_w_10_000_s_12_000 = 2.74e-11  mcrdlm4_cf_w_10_000_s_12_000 = 2.15e-11
+ mcrdlm4_ca_w_10_000_s_30_000 = 5.55e-06  mcrdlm4_cc_w_10_000_s_30_000 = 1.05e-11  mcrdlm4_cf_w_10_000_s_30_000 = 3.42e-11
+ mcrdlm4_ca_w_40_000_s_5_000 = 5.55e-06  mcrdlm4_cc_w_40_000_s_5_000 = 7.03e-11  mcrdlm4_cf_w_40_000_s_5_000 = 1.03e-11
+ mcrdlm4_ca_w_40_000_s_8_000 = 5.55e-06  mcrdlm4_cc_w_40_000_s_8_000 = 4.97e-11  mcrdlm4_cf_w_40_000_s_8_000 = 1.58e-11
+ mcrdlm4_ca_w_40_000_s_10_000 = 5.55e-06  mcrdlm4_cc_w_40_000_s_10_000 = 4.22e-11  mcrdlm4_cf_w_40_000_s_10_000 = 1.89e-11
+ mcrdlm4_ca_w_40_000_s_12_000 = 5.55e-06  mcrdlm4_cc_w_40_000_s_12_000 = 3.70e-11  mcrdlm4_cf_w_40_000_s_12_000 = 2.15e-11
+ mcrdlm4_ca_w_40_000_s_30_000 = 5.55e-06  mcrdlm4_cc_w_40_000_s_30_000 = 1.76e-11  mcrdlm4_cf_w_40_000_s_30_000 = 3.52e-11
+ mcrdlm5_ca_w_10_000_s_5_000 = 7.92e-06  mcrdlm5_cc_w_10_000_s_5_000 = 5.56e-11  mcrdlm5_cf_w_10_000_s_5_000 = 1.39e-11
+ mcrdlm5_ca_w_10_000_s_8_000 = 7.92e-06  mcrdlm5_cc_w_10_000_s_8_000 = 3.64e-11  mcrdlm5_cf_w_10_000_s_8_000 = 2.06e-11
+ mcrdlm5_ca_w_10_000_s_10_000 = 7.92e-06  mcrdlm5_cc_w_10_000_s_10_000 = 2.96e-11  mcrdlm5_cf_w_10_000_s_10_000 = 2.40e-11
+ mcrdlm5_ca_w_10_000_s_12_000 = 7.92e-06  mcrdlm5_cc_w_10_000_s_12_000 = 2.50e-11  mcrdlm5_cf_w_10_000_s_12_000 = 2.68e-11
+ mcrdlm5_ca_w_10_000_s_30_000 = 7.92e-06  mcrdlm5_cc_w_10_000_s_30_000 = 9.20e-12  mcrdlm5_cf_w_10_000_s_30_000 = 3.95e-11
+ mcrdlm5_ca_w_40_000_s_5_000 = 7.92e-06  mcrdlm5_cc_w_40_000_s_5_000 = 6.70e-11  mcrdlm5_cf_w_40_000_s_5_000 = 1.39e-11
+ mcrdlm5_ca_w_40_000_s_8_000 = 7.92e-06  mcrdlm5_cc_w_40_000_s_8_000 = 4.68e-11  mcrdlm5_cf_w_40_000_s_8_000 = 2.05e-11
+ mcrdlm5_ca_w_40_000_s_10_000 = 7.92e-06  mcrdlm5_cc_w_40_000_s_10_000 = 3.96e-11  mcrdlm5_cf_w_40_000_s_10_000 = 2.40e-11
+ mcrdlm5_ca_w_40_000_s_12_000 = 7.92e-06  mcrdlm5_cc_w_40_000_s_12_000 = 3.45e-11  mcrdlm5_cf_w_40_000_s_12_000 = 2.69e-11
+ mcrdlm5_ca_w_40_000_s_30_000 = 7.92e-06  mcrdlm5_cc_w_40_000_s_30_000 = 1.62e-11  mcrdlm5_cf_w_40_000_s_30_000 = 4.07e-11
+ mcl1p1f_ca_w_0_150_s_0_210 = 2.76e-04  mcl1p1f_cc_w_0_150_s_0_210 = 6.85e-11  mcl1p1f_cf_w_0_150_s_0_210 = 2.40e-11
+ mcl1p1f_ca_w_0_150_s_0_263 = 2.76e-04  mcl1p1f_cc_w_0_150_s_0_263 = 4.99e-11  mcl1p1f_cf_w_0_150_s_0_263 = 2.92e-11
+ mcl1p1f_ca_w_0_150_s_0_315 = 2.76e-04  mcl1p1f_cc_w_0_150_s_0_315 = 3.80e-11  mcl1p1f_cf_w_0_150_s_0_315 = 3.38e-11
+ mcl1p1f_ca_w_0_150_s_0_420 = 2.76e-04  mcl1p1f_cc_w_0_150_s_0_420 = 2.33e-11  mcl1p1f_cf_w_0_150_s_0_420 = 4.16e-11
+ mcl1p1f_ca_w_0_150_s_0_525 = 2.76e-04  mcl1p1f_cc_w_0_150_s_0_525 = 1.48e-11  mcl1p1f_cf_w_0_150_s_0_525 = 4.74e-11
+ mcl1p1f_ca_w_0_150_s_0_630 = 2.76e-04  mcl1p1f_cc_w_0_150_s_0_630 = 9.50e-12  mcl1p1f_cf_w_0_150_s_0_630 = 5.15e-11
+ mcl1p1f_ca_w_0_150_s_0_840 = 2.76e-04  mcl1p1f_cc_w_0_150_s_0_840 = 4.01e-12  mcl1p1f_cf_w_0_150_s_0_840 = 5.63e-11
+ mcl1p1f_ca_w_0_150_s_1_260 = 2.76e-04  mcl1p1f_cc_w_0_150_s_1_260 = 8.30e-13  mcl1p1f_cf_w_0_150_s_1_260 = 5.95e-11
+ mcl1p1f_ca_w_0_150_s_2_310 = 2.76e-04  mcl1p1f_cc_w_0_150_s_2_310 = 4.50e-14  mcl1p1f_cf_w_0_150_s_2_310 = 6.01e-11
+ mcl1p1f_ca_w_0_150_s_5_250 = 2.76e-04  mcl1p1f_cc_w_0_150_s_5_250 = 6.46e-27  mcl1p1f_cf_w_0_150_s_5_250 = 6.02e-11
+ mcl1p1f_ca_w_1_200_s_0_210 = 2.76e-04  mcl1p1f_cc_w_1_200_s_0_210 = 6.98e-11  mcl1p1f_cf_w_1_200_s_0_210 = 2.39e-11
+ mcl1p1f_ca_w_1_200_s_0_263 = 2.76e-04  mcl1p1f_cc_w_1_200_s_0_263 = 5.06e-11  mcl1p1f_cf_w_1_200_s_0_263 = 2.91e-11
+ mcl1p1f_ca_w_1_200_s_0_315 = 2.76e-04  mcl1p1f_cc_w_1_200_s_0_315 = 3.86e-11  mcl1p1f_cf_w_1_200_s_0_315 = 3.37e-11
+ mcl1p1f_ca_w_1_200_s_0_420 = 2.76e-04  mcl1p1f_cc_w_1_200_s_0_420 = 2.38e-11  mcl1p1f_cf_w_1_200_s_0_420 = 4.15e-11
+ mcl1p1f_ca_w_1_200_s_0_525 = 2.76e-04  mcl1p1f_cc_w_1_200_s_0_525 = 1.50e-11  mcl1p1f_cf_w_1_200_s_0_525 = 4.74e-11
+ mcl1p1f_ca_w_1_200_s_0_630 = 2.76e-04  mcl1p1f_cc_w_1_200_s_0_630 = 9.70e-12  mcl1p1f_cf_w_1_200_s_0_630 = 5.16e-11
+ mcl1p1f_ca_w_1_200_s_0_840 = 2.76e-04  mcl1p1f_cc_w_1_200_s_0_840 = 4.15e-12  mcl1p1f_cf_w_1_200_s_0_840 = 5.66e-11
+ mcl1p1f_ca_w_1_200_s_1_260 = 2.76e-04  mcl1p1f_cc_w_1_200_s_1_260 = 8.00e-13  mcl1p1f_cf_w_1_200_s_1_260 = 5.98e-11
+ mcl1p1f_ca_w_1_200_s_2_310 = 2.76e-04  mcl1p1f_cc_w_1_200_s_2_310 = 5.00e-14  mcl1p1f_cf_w_1_200_s_2_310 = 6.05e-11
+ mcl1p1f_ca_w_1_200_s_5_250 = 2.76e-04  mcl1p1f_cc_w_1_200_s_5_250 = 5.00e-14  mcl1p1f_cf_w_1_200_s_5_250 = 6.05e-11
+ mcm1p1f_ca_w_0_150_s_0_210 = 1.97e-04  mcm1p1f_cc_w_0_150_s_0_210 = 7.63e-11  mcm1p1f_cf_w_0_150_s_0_210 = 1.77e-11
+ mcm1p1f_ca_w_0_150_s_0_263 = 1.97e-04  mcm1p1f_cc_w_0_150_s_0_263 = 5.79e-11  mcm1p1f_cf_w_0_150_s_0_263 = 2.18e-11
+ mcm1p1f_ca_w_0_150_s_0_315 = 1.97e-04  mcm1p1f_cc_w_0_150_s_0_315 = 4.59e-11  mcm1p1f_cf_w_0_150_s_0_315 = 2.55e-11
+ mcm1p1f_ca_w_0_150_s_0_420 = 1.97e-04  mcm1p1f_cc_w_0_150_s_0_420 = 3.10e-11  mcm1p1f_cf_w_0_150_s_0_420 = 3.21e-11
+ mcm1p1f_ca_w_0_150_s_0_525 = 1.97e-04  mcm1p1f_cc_w_0_150_s_0_525 = 2.18e-11  mcm1p1f_cf_w_0_150_s_0_525 = 3.73e-11
+ mcm1p1f_ca_w_0_150_s_0_630 = 1.97e-04  mcm1p1f_cc_w_0_150_s_0_630 = 1.56e-11  mcm1p1f_cf_w_0_150_s_0_630 = 4.15e-11
+ mcm1p1f_ca_w_0_150_s_0_840 = 1.97e-04  mcm1p1f_cc_w_0_150_s_0_840 = 8.38e-12  mcm1p1f_cf_w_0_150_s_0_840 = 4.72e-11
+ mcm1p1f_ca_w_0_150_s_1_260 = 1.97e-04  mcm1p1f_cc_w_0_150_s_1_260 = 2.61e-12  mcm1p1f_cf_w_0_150_s_1_260 = 5.25e-11
+ mcm1p1f_ca_w_0_150_s_2_310 = 1.97e-04  mcm1p1f_cc_w_0_150_s_2_310 = 2.10e-13  mcm1p1f_cf_w_0_150_s_2_310 = 5.48e-11
+ mcm1p1f_ca_w_0_150_s_5_250 = 1.97e-04  mcm1p1f_cc_w_0_150_s_5_250 = 5.00e-15  mcm1p1f_cf_w_0_150_s_5_250 = 5.50e-11
+ mcm1p1f_ca_w_1_200_s_0_210 = 1.97e-04  mcm1p1f_cc_w_1_200_s_0_210 = 8.04e-11  mcm1p1f_cf_w_1_200_s_0_210 = 1.76e-11
+ mcm1p1f_ca_w_1_200_s_0_263 = 1.97e-04  mcm1p1f_cc_w_1_200_s_0_263 = 6.11e-11  mcm1p1f_cf_w_1_200_s_0_263 = 2.17e-11
+ mcm1p1f_ca_w_1_200_s_0_315 = 1.97e-04  mcm1p1f_cc_w_1_200_s_0_315 = 4.87e-11  mcm1p1f_cf_w_1_200_s_0_315 = 2.54e-11
+ mcm1p1f_ca_w_1_200_s_0_420 = 1.97e-04  mcm1p1f_cc_w_1_200_s_0_420 = 3.30e-11  mcm1p1f_cf_w_1_200_s_0_420 = 3.20e-11
+ mcm1p1f_ca_w_1_200_s_0_525 = 1.97e-04  mcm1p1f_cc_w_1_200_s_0_525 = 2.34e-11  mcm1p1f_cf_w_1_200_s_0_525 = 3.74e-11
+ mcm1p1f_ca_w_1_200_s_0_630 = 1.97e-04  mcm1p1f_cc_w_1_200_s_0_630 = 1.69e-11  mcm1p1f_cf_w_1_200_s_0_630 = 4.18e-11
+ mcm1p1f_ca_w_1_200_s_0_840 = 1.97e-04  mcm1p1f_cc_w_1_200_s_0_840 = 9.20e-12  mcm1p1f_cf_w_1_200_s_0_840 = 4.78e-11
+ mcm1p1f_ca_w_1_200_s_1_260 = 1.97e-04  mcm1p1f_cc_w_1_200_s_1_260 = 2.85e-12  mcm1p1f_cf_w_1_200_s_1_260 = 5.35e-11
+ mcm1p1f_ca_w_1_200_s_2_310 = 1.97e-04  mcm1p1f_cc_w_1_200_s_2_310 = 2.50e-13  mcm1p1f_cf_w_1_200_s_2_310 = 5.61e-11
+ mcm1p1f_ca_w_1_200_s_5_250 = 1.97e-04  mcm1p1f_cc_w_1_200_s_5_250 = 6.46e-27  mcm1p1f_cf_w_1_200_s_5_250 = 5.63e-11
+ mcm2p1f_ca_w_0_150_s_0_210 = 1.67e-04  mcm2p1f_cc_w_0_150_s_0_210 = 8.04e-11  mcm2p1f_cf_w_0_150_s_0_210 = 1.51e-11
+ mcm2p1f_ca_w_0_150_s_0_263 = 1.67e-04  mcm2p1f_cc_w_0_150_s_0_263 = 6.22e-11  mcm2p1f_cf_w_0_150_s_0_263 = 1.86e-11
+ mcm2p1f_ca_w_0_150_s_0_315 = 1.67e-04  mcm2p1f_cc_w_0_150_s_0_315 = 5.05e-11  mcm2p1f_cf_w_0_150_s_0_315 = 2.17e-11
+ mcm2p1f_ca_w_0_150_s_0_420 = 1.67e-04  mcm2p1f_cc_w_0_150_s_0_420 = 3.58e-11  mcm2p1f_cf_w_0_150_s_0_420 = 2.75e-11
+ mcm2p1f_ca_w_0_150_s_0_525 = 1.67e-04  mcm2p1f_cc_w_0_150_s_0_525 = 2.66e-11  mcm2p1f_cf_w_0_150_s_0_525 = 3.22e-11
+ mcm2p1f_ca_w_0_150_s_0_630 = 1.67e-04  mcm2p1f_cc_w_0_150_s_0_630 = 2.04e-11  mcm2p1f_cf_w_0_150_s_0_630 = 3.61e-11
+ mcm2p1f_ca_w_0_150_s_0_840 = 1.67e-04  mcm2p1f_cc_w_0_150_s_0_840 = 1.25e-11  mcm2p1f_cf_w_0_150_s_0_840 = 4.19e-11
+ mcm2p1f_ca_w_0_150_s_1_260 = 1.67e-04  mcm2p1f_cc_w_0_150_s_1_260 = 5.23e-12  mcm2p1f_cf_w_0_150_s_1_260 = 4.81e-11
+ mcm2p1f_ca_w_0_150_s_2_310 = 1.67e-04  mcm2p1f_cc_w_0_150_s_2_310 = 7.35e-13  mcm2p1f_cf_w_0_150_s_2_310 = 5.23e-11
+ mcm2p1f_ca_w_0_150_s_5_250 = 1.67e-04  mcm2p1f_cc_w_0_150_s_5_250 = 3.50e-14  mcm2p1f_cf_w_0_150_s_5_250 = 5.30e-11
+ mcm2p1f_ca_w_1_200_s_0_210 = 1.67e-04  mcm2p1f_cc_w_1_200_s_0_210 = 8.83e-11  mcm2p1f_cf_w_1_200_s_0_210 = 1.50e-11
+ mcm2p1f_ca_w_1_200_s_0_263 = 1.67e-04  mcm2p1f_cc_w_1_200_s_0_263 = 6.89e-11  mcm2p1f_cf_w_1_200_s_0_263 = 1.85e-11
+ mcm2p1f_ca_w_1_200_s_0_315 = 1.67e-04  mcm2p1f_cc_w_1_200_s_0_315 = 5.65e-11  mcm2p1f_cf_w_1_200_s_0_315 = 2.17e-11
+ mcm2p1f_ca_w_1_200_s_0_420 = 1.67e-04  mcm2p1f_cc_w_1_200_s_0_420 = 4.05e-11  mcm2p1f_cf_w_1_200_s_0_420 = 2.75e-11
+ mcm2p1f_ca_w_1_200_s_0_525 = 1.67e-04  mcm2p1f_cc_w_1_200_s_0_525 = 3.06e-11  mcm2p1f_cf_w_1_200_s_0_525 = 3.24e-11
+ mcm2p1f_ca_w_1_200_s_0_630 = 1.67e-04  mcm2p1f_cc_w_1_200_s_0_630 = 2.38e-11  mcm2p1f_cf_w_1_200_s_0_630 = 3.64e-11
+ mcm2p1f_ca_w_1_200_s_0_840 = 1.67e-04  mcm2p1f_cc_w_1_200_s_0_840 = 1.51e-11  mcm2p1f_cf_w_1_200_s_0_840 = 4.26e-11
+ mcm2p1f_ca_w_1_200_s_1_260 = 1.67e-04  mcm2p1f_cc_w_1_200_s_1_260 = 6.58e-12  mcm2p1f_cf_w_1_200_s_1_260 = 4.97e-11
+ mcm2p1f_ca_w_1_200_s_2_310 = 1.67e-04  mcm2p1f_cc_w_1_200_s_2_310 = 9.70e-13  mcm2p1f_cf_w_1_200_s_2_310 = 5.50e-11
+ mcm2p1f_ca_w_1_200_s_5_250 = 1.67e-04  mcm2p1f_cc_w_1_200_s_5_250 = 5.00e-15  mcm2p1f_cf_w_1_200_s_5_250 = 5.59e-11
+ mcm3p1f_ca_w_0_150_s_0_210 = 1.55e-04  mcm3p1f_cc_w_0_150_s_0_210 = 8.21e-11  mcm3p1f_cf_w_0_150_s_0_210 = 1.40e-11
+ mcm3p1f_ca_w_0_150_s_0_263 = 1.55e-04  mcm3p1f_cc_w_0_150_s_0_263 = 6.42e-11  mcm3p1f_cf_w_0_150_s_0_263 = 1.72e-11
+ mcm3p1f_ca_w_0_150_s_0_315 = 1.55e-04  mcm3p1f_cc_w_0_150_s_0_315 = 5.26e-11  mcm3p1f_cf_w_0_150_s_0_315 = 2.01e-11
+ mcm3p1f_ca_w_0_150_s_0_420 = 1.55e-04  mcm3p1f_cc_w_0_150_s_0_420 = 3.81e-11  mcm3p1f_cf_w_0_150_s_0_420 = 2.55e-11
+ mcm3p1f_ca_w_0_150_s_0_525 = 1.55e-04  mcm3p1f_cc_w_0_150_s_0_525 = 2.92e-11  mcm3p1f_cf_w_0_150_s_0_525 = 3.00e-11
+ mcm3p1f_ca_w_0_150_s_0_630 = 1.55e-04  mcm3p1f_cc_w_0_150_s_0_630 = 2.30e-11  mcm3p1f_cf_w_0_150_s_0_630 = 3.36e-11
+ mcm3p1f_ca_w_0_150_s_0_840 = 1.55e-04  mcm3p1f_cc_w_0_150_s_0_840 = 1.50e-11  mcm3p1f_cf_w_0_150_s_0_840 = 3.93e-11
+ mcm3p1f_ca_w_0_150_s_1_260 = 1.55e-04  mcm3p1f_cc_w_0_150_s_1_260 = 7.16e-12  mcm3p1f_cf_w_0_150_s_1_260 = 4.59e-11
+ mcm3p1f_ca_w_0_150_s_2_310 = 1.55e-04  mcm3p1f_cc_w_0_150_s_2_310 = 1.51e-12  mcm3p1f_cf_w_0_150_s_2_310 = 5.10e-11
+ mcm3p1f_ca_w_0_150_s_5_250 = 1.55e-04  mcm3p1f_cc_w_0_150_s_5_250 = 3.00e-14  mcm3p1f_cf_w_0_150_s_5_250 = 5.24e-11
+ mcm3p1f_ca_w_1_200_s_0_210 = 1.55e-04  mcm3p1f_cc_w_1_200_s_0_210 = 9.30e-11  mcm3p1f_cf_w_1_200_s_0_210 = 1.39e-11
+ mcm3p1f_ca_w_1_200_s_0_263 = 1.55e-04  mcm3p1f_cc_w_1_200_s_0_263 = 7.37e-11  mcm3p1f_cf_w_1_200_s_0_263 = 1.72e-11
+ mcm3p1f_ca_w_1_200_s_0_315 = 1.55e-04  mcm3p1f_cc_w_1_200_s_0_315 = 6.13e-11  mcm3p1f_cf_w_1_200_s_0_315 = 2.01e-11
+ mcm3p1f_ca_w_1_200_s_0_420 = 1.55e-04  mcm3p1f_cc_w_1_200_s_0_420 = 4.53e-11  mcm3p1f_cf_w_1_200_s_0_420 = 2.55e-11
+ mcm3p1f_ca_w_1_200_s_0_525 = 1.55e-04  mcm3p1f_cc_w_1_200_s_0_525 = 3.54e-11  mcm3p1f_cf_w_1_200_s_0_525 = 3.00e-11
+ mcm3p1f_ca_w_1_200_s_0_630 = 1.55e-04  mcm3p1f_cc_w_1_200_s_0_630 = 2.84e-11  mcm3p1f_cf_w_1_200_s_0_630 = 3.39e-11
+ mcm3p1f_ca_w_1_200_s_0_840 = 1.55e-04  mcm3p1f_cc_w_1_200_s_0_840 = 1.93e-11  mcm3p1f_cf_w_1_200_s_0_840 = 4.00e-11
+ mcm3p1f_ca_w_1_200_s_1_260 = 1.55e-04  mcm3p1f_cc_w_1_200_s_1_260 = 9.89e-12  mcm3p1f_cf_w_1_200_s_1_260 = 4.74e-11
+ mcm3p1f_ca_w_1_200_s_2_310 = 1.55e-04  mcm3p1f_cc_w_1_200_s_2_310 = 2.29e-12  mcm3p1f_cf_w_1_200_s_2_310 = 5.44e-11
+ mcm3p1f_ca_w_1_200_s_5_250 = 1.55e-04  mcm3p1f_cc_w_1_200_s_5_250 = 1.00e-13  mcm3p1f_cf_w_1_200_s_5_250 = 5.66e-11
+ mcm4p1f_ca_w_0_150_s_0_210 = 1.48e-04  mcm4p1f_cc_w_0_150_s_0_210 = 8.32e-11  mcm4p1f_cf_w_0_150_s_0_210 = 1.33e-11
+ mcm4p1f_ca_w_0_150_s_0_263 = 1.48e-04  mcm4p1f_cc_w_0_150_s_0_263 = 6.54e-11  mcm4p1f_cf_w_0_150_s_0_263 = 1.63e-11
+ mcm4p1f_ca_w_0_150_s_0_315 = 1.48e-04  mcm4p1f_cc_w_0_150_s_0_315 = 5.41e-11  mcm4p1f_cf_w_0_150_s_0_315 = 1.91e-11
+ mcm4p1f_ca_w_0_150_s_0_420 = 1.48e-04  mcm4p1f_cc_w_0_150_s_0_420 = 3.97e-11  mcm4p1f_cf_w_0_150_s_0_420 = 2.42e-11
+ mcm4p1f_ca_w_0_150_s_0_525 = 1.48e-04  mcm4p1f_cc_w_0_150_s_0_525 = 3.10e-11  mcm4p1f_cf_w_0_150_s_0_525 = 2.84e-11
+ mcm4p1f_ca_w_0_150_s_0_630 = 1.48e-04  mcm4p1f_cc_w_0_150_s_0_630 = 2.49e-11  mcm4p1f_cf_w_0_150_s_0_630 = 3.19e-11
+ mcm4p1f_ca_w_0_150_s_0_840 = 1.48e-04  mcm4p1f_cc_w_0_150_s_0_840 = 1.70e-11  mcm4p1f_cf_w_0_150_s_0_840 = 3.75e-11
+ mcm4p1f_ca_w_0_150_s_1_260 = 1.48e-04  mcm4p1f_cc_w_0_150_s_1_260 = 8.72e-12  mcm4p1f_cf_w_0_150_s_1_260 = 4.43e-11
+ mcm4p1f_ca_w_0_150_s_2_310 = 1.48e-04  mcm4p1f_cc_w_0_150_s_2_310 = 2.41e-12  mcm4p1f_cf_w_0_150_s_2_310 = 4.99e-11
+ mcm4p1f_ca_w_0_150_s_5_250 = 1.48e-04  mcm4p1f_cc_w_0_150_s_5_250 = 1.70e-13  mcm4p1f_cf_w_0_150_s_5_250 = 5.21e-11
+ mcm4p1f_ca_w_1_200_s_0_210 = 1.48e-04  mcm4p1f_cc_w_1_200_s_0_210 = 9.68e-11  mcm4p1f_cf_w_1_200_s_0_210 = 1.33e-11
+ mcm4p1f_ca_w_1_200_s_0_263 = 1.48e-04  mcm4p1f_cc_w_1_200_s_0_263 = 7.75e-11  mcm4p1f_cf_w_1_200_s_0_263 = 1.63e-11
+ mcm4p1f_ca_w_1_200_s_0_315 = 1.48e-04  mcm4p1f_cc_w_1_200_s_0_315 = 6.51e-11  mcm4p1f_cf_w_1_200_s_0_315 = 1.91e-11
+ mcm4p1f_ca_w_1_200_s_0_420 = 1.48e-04  mcm4p1f_cc_w_1_200_s_0_420 = 4.92e-11  mcm4p1f_cf_w_1_200_s_0_420 = 2.41e-11
+ mcm4p1f_ca_w_1_200_s_0_525 = 1.48e-04  mcm4p1f_cc_w_1_200_s_0_525 = 3.94e-11  mcm4p1f_cf_w_1_200_s_0_525 = 2.85e-11
+ mcm4p1f_ca_w_1_200_s_0_630 = 1.48e-04  mcm4p1f_cc_w_1_200_s_0_630 = 3.24e-11  mcm4p1f_cf_w_1_200_s_0_630 = 3.22e-11
+ mcm4p1f_ca_w_1_200_s_0_840 = 1.48e-04  mcm4p1f_cc_w_1_200_s_0_840 = 2.32e-11  mcm4p1f_cf_w_1_200_s_0_840 = 3.81e-11
+ mcm4p1f_ca_w_1_200_s_1_260 = 1.48e-04  mcm4p1f_cc_w_1_200_s_1_260 = 1.32e-11  mcm4p1f_cf_w_1_200_s_1_260 = 4.58e-11
+ mcm4p1f_ca_w_1_200_s_2_310 = 1.48e-04  mcm4p1f_cc_w_1_200_s_2_310 = 4.16e-12  mcm4p1f_cf_w_1_200_s_2_310 = 5.38e-11
+ mcm4p1f_ca_w_1_200_s_5_250 = 1.48e-04  mcm4p1f_cc_w_1_200_s_5_250 = 2.85e-13  mcm4p1f_cf_w_1_200_s_5_250 = 5.76e-11
+ mcm5p1f_ca_w_0_150_s_0_210 = 1.44e-04  mcm5p1f_cc_w_0_150_s_0_210 = 8.37e-11  mcm5p1f_cf_w_0_150_s_0_210 = 1.30e-11
+ mcm5p1f_ca_w_0_150_s_0_263 = 1.44e-04  mcm5p1f_cc_w_0_150_s_0_263 = 6.59e-11  mcm5p1f_cf_w_0_150_s_0_263 = 1.59e-11
+ mcm5p1f_ca_w_0_150_s_0_315 = 1.44e-04  mcm5p1f_cc_w_0_150_s_0_315 = 5.47e-11  mcm5p1f_cf_w_0_150_s_0_315 = 1.86e-11
+ mcm5p1f_ca_w_0_150_s_0_420 = 1.44e-04  mcm5p1f_cc_w_0_150_s_0_420 = 4.04e-11  mcm5p1f_cf_w_0_150_s_0_420 = 2.36e-11
+ mcm5p1f_ca_w_0_150_s_0_525 = 1.44e-04  mcm5p1f_cc_w_0_150_s_0_525 = 3.18e-11  mcm5p1f_cf_w_0_150_s_0_525 = 2.77e-11
+ mcm5p1f_ca_w_0_150_s_0_630 = 1.44e-04  mcm5p1f_cc_w_0_150_s_0_630 = 2.58e-11  mcm5p1f_cf_w_0_150_s_0_630 = 3.11e-11
+ mcm5p1f_ca_w_0_150_s_0_840 = 1.44e-04  mcm5p1f_cc_w_0_150_s_0_840 = 1.79e-11  mcm5p1f_cf_w_0_150_s_0_840 = 3.66e-11
+ mcm5p1f_ca_w_0_150_s_1_260 = 1.44e-04  mcm5p1f_cc_w_0_150_s_1_260 = 9.51e-12  mcm5p1f_cf_w_0_150_s_1_260 = 4.35e-11
+ mcm5p1f_ca_w_0_150_s_2_310 = 1.44e-04  mcm5p1f_cc_w_0_150_s_2_310 = 3.02e-12  mcm5p1f_cf_w_0_150_s_2_310 = 4.93e-11
+ mcm5p1f_ca_w_0_150_s_5_250 = 1.44e-04  mcm5p1f_cc_w_0_150_s_5_250 = 3.19e-13  mcm5p1f_cf_w_0_150_s_5_250 = 5.20e-11
+ mcm5p1f_ca_w_1_200_s_0_210 = 1.44e-04  mcm5p1f_cc_w_1_200_s_0_210 = 9.86e-11  mcm5p1f_cf_w_1_200_s_0_210 = 1.29e-11
+ mcm5p1f_ca_w_1_200_s_0_263 = 1.44e-04  mcm5p1f_cc_w_1_200_s_0_263 = 7.95e-11  mcm5p1f_cf_w_1_200_s_0_263 = 1.59e-11
+ mcm5p1f_ca_w_1_200_s_0_315 = 1.44e-04  mcm5p1f_cc_w_1_200_s_0_315 = 6.71e-11  mcm5p1f_cf_w_1_200_s_0_315 = 1.86e-11
+ mcm5p1f_ca_w_1_200_s_0_420 = 1.44e-04  mcm5p1f_cc_w_1_200_s_0_420 = 5.14e-11  mcm5p1f_cf_w_1_200_s_0_420 = 2.35e-11
+ mcm5p1f_ca_w_1_200_s_0_525 = 1.44e-04  mcm5p1f_cc_w_1_200_s_0_525 = 4.16e-11  mcm5p1f_cf_w_1_200_s_0_525 = 2.77e-11
+ mcm5p1f_ca_w_1_200_s_0_630 = 1.44e-04  mcm5p1f_cc_w_1_200_s_0_630 = 3.46e-11  mcm5p1f_cf_w_1_200_s_0_630 = 3.14e-11
+ mcm5p1f_ca_w_1_200_s_0_840 = 1.44e-04  mcm5p1f_cc_w_1_200_s_0_840 = 2.53e-11  mcm5p1f_cf_w_1_200_s_0_840 = 3.72e-11
+ mcm5p1f_ca_w_1_200_s_1_260 = 1.44e-04  mcm5p1f_cc_w_1_200_s_1_260 = 1.52e-11  mcm5p1f_cf_w_1_200_s_1_260 = 4.48e-11
+ mcm5p1f_ca_w_1_200_s_2_310 = 1.44e-04  mcm5p1f_cc_w_1_200_s_2_310 = 5.53e-12  mcm5p1f_cf_w_1_200_s_2_310 = 5.34e-11
+ mcm5p1f_ca_w_1_200_s_5_250 = 1.44e-04  mcm5p1f_cc_w_1_200_s_5_250 = 6.50e-13  mcm5p1f_cf_w_1_200_s_5_250 = 5.81e-11
+ mcrdlp1f_ca_w_0_150_s_0_210 = 1.39e-04  mcrdlp1f_cc_w_0_150_s_0_210 = 8.44e-11  mcrdlp1f_cf_w_0_150_s_0_210 = 1.25e-11
+ mcrdlp1f_ca_w_0_150_s_0_263 = 1.39e-04  mcrdlp1f_cc_w_0_150_s_0_263 = 6.67e-11  mcrdlp1f_cf_w_0_150_s_0_263 = 1.53e-11
+ mcrdlp1f_ca_w_0_150_s_0_315 = 1.39e-04  mcrdlp1f_cc_w_0_150_s_0_315 = 5.56e-11  mcrdlp1f_cf_w_0_150_s_0_315 = 1.79e-11
+ mcrdlp1f_ca_w_0_150_s_0_420 = 1.39e-04  mcrdlp1f_cc_w_0_150_s_0_420 = 4.14e-11  mcrdlp1f_cf_w_0_150_s_0_420 = 2.27e-11
+ mcrdlp1f_ca_w_0_150_s_0_525 = 1.39e-04  mcrdlp1f_cc_w_0_150_s_0_525 = 3.30e-11  mcrdlp1f_cf_w_0_150_s_0_525 = 2.66e-11
+ mcrdlp1f_ca_w_0_150_s_0_630 = 1.39e-04  mcrdlp1f_cc_w_0_150_s_0_630 = 2.72e-11  mcrdlp1f_cf_w_0_150_s_0_630 = 3.00e-11
+ mcrdlp1f_ca_w_0_150_s_0_840 = 1.39e-04  mcrdlp1f_cc_w_0_150_s_0_840 = 1.93e-11  mcrdlp1f_cf_w_0_150_s_0_840 = 3.53e-11
+ mcrdlp1f_ca_w_0_150_s_1_260 = 1.39e-04  mcrdlp1f_cc_w_0_150_s_1_260 = 1.07e-11  mcrdlp1f_cf_w_0_150_s_1_260 = 4.24e-11
+ mcrdlp1f_ca_w_0_150_s_2_310 = 1.39e-04  mcrdlp1f_cc_w_0_150_s_2_310 = 4.08e-12  mcrdlp1f_cf_w_0_150_s_2_310 = 4.84e-11
+ mcrdlp1f_ca_w_0_150_s_5_250 = 1.39e-04  mcrdlp1f_cc_w_0_150_s_5_250 = 7.44e-13  mcrdlp1f_cf_w_0_150_s_5_250 = 5.17e-11
+ mcrdlp1f_ca_w_1_200_s_0_210 = 1.39e-04  mcrdlp1f_cc_w_1_200_s_0_210 = 1.01e-10  mcrdlp1f_cf_w_1_200_s_0_210 = 1.24e-11
+ mcrdlp1f_ca_w_1_200_s_0_263 = 1.39e-04  mcrdlp1f_cc_w_1_200_s_0_263 = 8.24e-11  mcrdlp1f_cf_w_1_200_s_0_263 = 1.53e-11
+ mcrdlp1f_ca_w_1_200_s_0_315 = 1.39e-04  mcrdlp1f_cc_w_1_200_s_0_315 = 7.02e-11  mcrdlp1f_cf_w_1_200_s_0_315 = 1.79e-11
+ mcrdlp1f_ca_w_1_200_s_0_420 = 1.39e-04  mcrdlp1f_cc_w_1_200_s_0_420 = 5.45e-11  mcrdlp1f_cf_w_1_200_s_0_420 = 2.26e-11
+ mcrdlp1f_ca_w_1_200_s_0_525 = 1.39e-04  mcrdlp1f_cc_w_1_200_s_0_525 = 4.48e-11  mcrdlp1f_cf_w_1_200_s_0_525 = 2.67e-11
+ mcrdlp1f_ca_w_1_200_s_0_630 = 1.39e-04  mcrdlp1f_cc_w_1_200_s_0_630 = 3.79e-11  mcrdlp1f_cf_w_1_200_s_0_630 = 3.02e-11
+ mcrdlp1f_ca_w_1_200_s_0_840 = 1.39e-04  mcrdlp1f_cc_w_1_200_s_0_840 = 2.88e-11  mcrdlp1f_cf_w_1_200_s_0_840 = 3.59e-11
+ mcrdlp1f_ca_w_1_200_s_1_260 = 1.39e-04  mcrdlp1f_cc_w_1_200_s_1_260 = 1.86e-11  mcrdlp1f_cf_w_1_200_s_1_260 = 4.35e-11
+ mcrdlp1f_ca_w_1_200_s_2_310 = 1.39e-04  mcrdlp1f_cc_w_1_200_s_2_310 = 8.14e-12  mcrdlp1f_cf_w_1_200_s_2_310 = 5.27e-11
+ mcrdlp1f_ca_w_1_200_s_5_250 = 1.39e-04  mcrdlp1f_cc_w_1_200_s_5_250 = 1.81e-12  mcrdlp1f_cf_w_1_200_s_5_250 = 5.88e-11
+ mcm1l1f_ca_w_0_170_s_0_180 = 2.08e-04  mcm1l1f_cc_w_0_170_s_0_180 = 7.61e-11  mcm1l1f_cf_w_0_170_s_0_180 = 1.49e-11
+ mcm1l1f_ca_w_0_170_s_0_225 = 2.08e-04  mcm1l1f_cc_w_0_170_s_0_225 = 5.90e-11  mcm1l1f_cf_w_0_170_s_0_225 = 1.86e-11
+ mcm1l1f_ca_w_0_170_s_0_270 = 2.08e-04  mcm1l1f_cc_w_0_170_s_0_270 = 4.78e-11  mcm1l1f_cf_w_0_170_s_0_270 = 2.19e-11
+ mcm1l1f_ca_w_0_170_s_0_360 = 2.08e-04  mcm1l1f_cc_w_0_170_s_0_360 = 3.32e-11  mcm1l1f_cf_w_0_170_s_0_360 = 2.79e-11
+ mcm1l1f_ca_w_0_170_s_0_450 = 2.08e-04  mcm1l1f_cc_w_0_170_s_0_450 = 2.42e-11  mcm1l1f_cf_w_0_170_s_0_450 = 3.28e-11
+ mcm1l1f_ca_w_0_170_s_0_540 = 2.08e-04  mcm1l1f_cc_w_0_170_s_0_540 = 1.81e-11  mcm1l1f_cf_w_0_170_s_0_540 = 3.70e-11
+ mcm1l1f_ca_w_0_170_s_0_720 = 2.08e-04  mcm1l1f_cc_w_0_170_s_0_720 = 1.04e-11  mcm1l1f_cf_w_0_170_s_0_720 = 4.28e-11
+ mcm1l1f_ca_w_0_170_s_1_080 = 2.08e-04  mcm1l1f_cc_w_0_170_s_1_080 = 3.69e-12  mcm1l1f_cf_w_0_170_s_1_080 = 4.87e-11
+ mcm1l1f_ca_w_0_170_s_1_980 = 2.08e-04  mcm1l1f_cc_w_0_170_s_1_980 = 3.80e-13  mcm1l1f_cf_w_0_170_s_1_980 = 5.19e-11
+ mcm1l1f_ca_w_0_170_s_4_500 = 2.08e-04  mcm1l1f_cc_w_0_170_s_4_500 = 3.50e-14  mcm1l1f_cf_w_0_170_s_4_500 = 5.23e-11
+ mcm1l1f_ca_w_1_360_s_0_180 = 2.08e-04  mcm1l1f_cc_w_1_360_s_0_180 = 7.97e-11  mcm1l1f_cf_w_1_360_s_0_180 = 1.48e-11
+ mcm1l1f_ca_w_1_360_s_0_225 = 2.08e-04  mcm1l1f_cc_w_1_360_s_0_225 = 6.23e-11  mcm1l1f_cf_w_1_360_s_0_225 = 1.85e-11
+ mcm1l1f_ca_w_1_360_s_0_270 = 2.08e-04  mcm1l1f_cc_w_1_360_s_0_270 = 5.05e-11  mcm1l1f_cf_w_1_360_s_0_270 = 2.18e-11
+ mcm1l1f_ca_w_1_360_s_0_360 = 2.08e-04  mcm1l1f_cc_w_1_360_s_0_360 = 3.55e-11  mcm1l1f_cf_w_1_360_s_0_360 = 2.79e-11
+ mcm1l1f_ca_w_1_360_s_0_450 = 2.08e-04  mcm1l1f_cc_w_1_360_s_0_450 = 2.61e-11  mcm1l1f_cf_w_1_360_s_0_450 = 3.29e-11
+ mcm1l1f_ca_w_1_360_s_0_540 = 2.08e-04  mcm1l1f_cc_w_1_360_s_0_540 = 1.96e-11  mcm1l1f_cf_w_1_360_s_0_540 = 3.71e-11
+ mcm1l1f_ca_w_1_360_s_0_720 = 2.08e-04  mcm1l1f_cc_w_1_360_s_0_720 = 1.14e-11  mcm1l1f_cf_w_1_360_s_0_720 = 4.31e-11
+ mcm1l1f_ca_w_1_360_s_1_080 = 2.08e-04  mcm1l1f_cc_w_1_360_s_1_080 = 4.16e-12  mcm1l1f_cf_w_1_360_s_1_080 = 4.95e-11
+ mcm1l1f_ca_w_1_360_s_1_980 = 2.08e-04  mcm1l1f_cc_w_1_360_s_1_980 = 4.20e-13  mcm1l1f_cf_w_1_360_s_1_980 = 5.31e-11
+ mcm1l1f_ca_w_1_360_s_4_500 = 2.08e-04  mcm1l1f_cc_w_1_360_s_4_500 = 2.00e-14  mcm1l1f_cf_w_1_360_s_4_500 = 5.34e-11
+ mcm1l1d_ca_w_0_170_s_0_180 = 2.29e-04  mcm1l1d_cc_w_0_170_s_0_180 = 7.36e-11  mcm1l1d_cf_w_0_170_s_0_180 = 1.65e-11
+ mcm1l1d_ca_w_0_170_s_0_225 = 2.29e-04  mcm1l1d_cc_w_0_170_s_0_225 = 5.64e-11  mcm1l1d_cf_w_0_170_s_0_225 = 2.04e-11
+ mcm1l1d_ca_w_0_170_s_0_270 = 2.29e-04  mcm1l1d_cc_w_0_170_s_0_270 = 4.50e-11  mcm1l1d_cf_w_0_170_s_0_270 = 2.41e-11
+ mcm1l1d_ca_w_0_170_s_0_360 = 2.29e-04  mcm1l1d_cc_w_0_170_s_0_360 = 3.04e-11  mcm1l1d_cf_w_0_170_s_0_360 = 3.06e-11
+ mcm1l1d_ca_w_0_170_s_0_450 = 2.29e-04  mcm1l1d_cc_w_0_170_s_0_450 = 2.14e-11  mcm1l1d_cf_w_0_170_s_0_450 = 3.58e-11
+ mcm1l1d_ca_w_0_170_s_0_540 = 2.29e-04  mcm1l1d_cc_w_0_170_s_0_540 = 1.55e-11  mcm1l1d_cf_w_0_170_s_0_540 = 4.00e-11
+ mcm1l1d_ca_w_0_170_s_0_720 = 2.29e-04  mcm1l1d_cc_w_0_170_s_0_720 = 8.23e-12  mcm1l1d_cf_w_0_170_s_0_720 = 4.58e-11
+ mcm1l1d_ca_w_0_170_s_1_080 = 2.29e-04  mcm1l1d_cc_w_0_170_s_1_080 = 2.46e-12  mcm1l1d_cf_w_0_170_s_1_080 = 5.11e-11
+ mcm1l1d_ca_w_0_170_s_1_980 = 2.29e-04  mcm1l1d_cc_w_0_170_s_1_980 = 2.00e-13  mcm1l1d_cf_w_0_170_s_1_980 = 5.33e-11
+ mcm1l1d_ca_w_0_170_s_4_500 = 2.29e-04  mcm1l1d_cc_w_0_170_s_4_500 = 0.00e+00  mcm1l1d_cf_w_0_170_s_4_500 = 5.34e-11
+ mcm1l1d_ca_w_1_360_s_0_180 = 2.29e-04  mcm1l1d_cc_w_1_360_s_0_180 = 7.63e-11  mcm1l1d_cf_w_1_360_s_0_180 = 1.63e-11
+ mcm1l1d_ca_w_1_360_s_0_225 = 2.29e-04  mcm1l1d_cc_w_1_360_s_0_225 = 5.86e-11  mcm1l1d_cf_w_1_360_s_0_225 = 2.03e-11
+ mcm1l1d_ca_w_1_360_s_0_270 = 2.29e-04  mcm1l1d_cc_w_1_360_s_0_270 = 4.68e-11  mcm1l1d_cf_w_1_360_s_0_270 = 2.40e-11
+ mcm1l1d_ca_w_1_360_s_0_360 = 2.29e-04  mcm1l1d_cc_w_1_360_s_0_360 = 3.17e-11  mcm1l1d_cf_w_1_360_s_0_360 = 3.05e-11
+ mcm1l1d_ca_w_1_360_s_0_450 = 2.29e-04  mcm1l1d_cc_w_1_360_s_0_450 = 2.25e-11  mcm1l1d_cf_w_1_360_s_0_450 = 3.57e-11
+ mcm1l1d_ca_w_1_360_s_0_540 = 2.29e-04  mcm1l1d_cc_w_1_360_s_0_540 = 1.62e-11  mcm1l1d_cf_w_1_360_s_0_540 = 4.00e-11
+ mcm1l1d_ca_w_1_360_s_0_720 = 2.29e-04  mcm1l1d_cc_w_1_360_s_0_720 = 8.70e-12  mcm1l1d_cf_w_1_360_s_0_720 = 4.60e-11
+ mcm1l1d_ca_w_1_360_s_1_080 = 2.29e-04  mcm1l1d_cc_w_1_360_s_1_080 = 2.60e-12  mcm1l1d_cf_w_1_360_s_1_080 = 5.15e-11
+ mcm1l1d_ca_w_1_360_s_1_980 = 2.29e-04  mcm1l1d_cc_w_1_360_s_1_980 = 2.00e-13  mcm1l1d_cf_w_1_360_s_1_980 = 5.39e-11
+ mcm1l1d_ca_w_1_360_s_4_500 = 2.29e-04  mcm1l1d_cc_w_1_360_s_4_500 = 0.00e+00  mcm1l1d_cf_w_1_360_s_4_500 = 5.40e-11
+ mcm1l1p1_ca_w_0_170_s_0_180 = 3.04e-04  mcm1l1p1_cc_w_0_170_s_0_180 = 6.69e-11  mcm1l1p1_cf_w_0_170_s_0_180 = 2.16e-11
+ mcm1l1p1_ca_w_0_170_s_0_225 = 3.04e-04  mcm1l1p1_cc_w_0_170_s_0_225 = 4.96e-11  mcm1l1p1_cf_w_0_170_s_0_225 = 2.67e-11
+ mcm1l1p1_ca_w_0_170_s_0_270 = 3.04e-04  mcm1l1p1_cc_w_0_170_s_0_270 = 3.82e-11  mcm1l1p1_cf_w_0_170_s_0_270 = 3.13e-11
+ mcm1l1p1_ca_w_0_170_s_0_360 = 3.04e-04  mcm1l1p1_cc_w_0_170_s_0_360 = 2.40e-11  mcm1l1p1_cf_w_0_170_s_0_360 = 3.92e-11
+ mcm1l1p1_ca_w_0_170_s_0_450 = 3.04e-04  mcm1l1p1_cc_w_0_170_s_0_450 = 1.55e-11  mcm1l1p1_cf_w_0_170_s_0_450 = 4.49e-11
+ mcm1l1p1_ca_w_0_170_s_0_540 = 3.04e-04  mcm1l1p1_cc_w_0_170_s_0_540 = 1.02e-11  mcm1l1p1_cf_w_0_170_s_0_540 = 4.92e-11
+ mcm1l1p1_ca_w_0_170_s_0_720 = 3.04e-04  mcm1l1p1_cc_w_0_170_s_0_720 = 4.44e-12  mcm1l1p1_cf_w_0_170_s_0_720 = 5.42e-11
+ mcm1l1p1_ca_w_0_170_s_1_080 = 3.04e-04  mcm1l1p1_cc_w_0_170_s_1_080 = 8.85e-13  mcm1l1p1_cf_w_0_170_s_1_080 = 5.76e-11
+ mcm1l1p1_ca_w_0_170_s_1_980 = 3.04e-04  mcm1l1p1_cc_w_0_170_s_1_980 = 5.50e-14  mcm1l1p1_cf_w_0_170_s_1_980 = 5.85e-11
+ mcm1l1p1_ca_w_0_170_s_4_500 = 3.04e-04  mcm1l1p1_cc_w_0_170_s_4_500 = 5.00e-15  mcm1l1p1_cf_w_0_170_s_4_500 = 5.85e-11
+ mcm1l1p1_ca_w_1_360_s_0_180 = 3.04e-04  mcm1l1p1_cc_w_1_360_s_0_180 = 6.76e-11  mcm1l1p1_cf_w_1_360_s_0_180 = 2.13e-11
+ mcm1l1p1_ca_w_1_360_s_0_225 = 3.04e-04  mcm1l1p1_cc_w_1_360_s_0_225 = 5.01e-11  mcm1l1p1_cf_w_1_360_s_0_225 = 2.64e-11
+ mcm1l1p1_ca_w_1_360_s_0_270 = 3.04e-04  mcm1l1p1_cc_w_1_360_s_0_270 = 3.88e-11  mcm1l1p1_cf_w_1_360_s_0_270 = 3.10e-11
+ mcm1l1p1_ca_w_1_360_s_0_360 = 3.04e-04  mcm1l1p1_cc_w_1_360_s_0_360 = 2.43e-11  mcm1l1p1_cf_w_1_360_s_0_360 = 3.88e-11
+ mcm1l1p1_ca_w_1_360_s_0_450 = 3.04e-04  mcm1l1p1_cc_w_1_360_s_0_450 = 1.58e-11  mcm1l1p1_cf_w_1_360_s_0_450 = 4.47e-11
+ mcm1l1p1_ca_w_1_360_s_0_540 = 3.04e-04  mcm1l1p1_cc_w_1_360_s_0_540 = 1.04e-11  mcm1l1p1_cf_w_1_360_s_0_540 = 4.90e-11
+ mcm1l1p1_ca_w_1_360_s_0_720 = 3.04e-04  mcm1l1p1_cc_w_1_360_s_0_720 = 4.55e-12  mcm1l1p1_cf_w_1_360_s_0_720 = 5.40e-11
+ mcm1l1p1_ca_w_1_360_s_1_080 = 3.04e-04  mcm1l1p1_cc_w_1_360_s_1_080 = 9.00e-13  mcm1l1p1_cf_w_1_360_s_1_080 = 5.75e-11
+ mcm1l1p1_ca_w_1_360_s_1_980 = 3.04e-04  mcm1l1p1_cc_w_1_360_s_1_980 = 5.00e-14  mcm1l1p1_cf_w_1_360_s_1_980 = 5.84e-11
+ mcm1l1p1_ca_w_1_360_s_4_500 = 3.04e-04  mcm1l1p1_cc_w_1_360_s_4_500 = 2.58e-26  mcm1l1p1_cf_w_1_360_s_4_500 = 5.83e-11
+ mcm2l1f_ca_w_0_170_s_0_180 = 9.12e-05  mcm2l1f_cc_w_0_170_s_0_180 = 8.69e-11  mcm2l1f_cf_w_0_170_s_0_180 = 6.94e-12
+ mcm2l1f_ca_w_0_170_s_0_225 = 9.12e-05  mcm2l1f_cc_w_0_170_s_0_225 = 7.04e-11  mcm2l1f_cf_w_0_170_s_0_225 = 8.82e-12
+ mcm2l1f_ca_w_0_170_s_0_270 = 9.12e-05  mcm2l1f_cc_w_0_170_s_0_270 = 5.92e-11  mcm2l1f_cf_w_0_170_s_0_270 = 1.06e-11
+ mcm2l1f_ca_w_0_170_s_0_360 = 9.12e-05  mcm2l1f_cc_w_0_170_s_0_360 = 4.47e-11  mcm2l1f_cf_w_0_170_s_0_360 = 1.42e-11
+ mcm2l1f_ca_w_0_170_s_0_450 = 9.12e-05  mcm2l1f_cc_w_0_170_s_0_450 = 3.54e-11  mcm2l1f_cf_w_0_170_s_0_450 = 1.74e-11
+ mcm2l1f_ca_w_0_170_s_0_540 = 9.12e-05  mcm2l1f_cc_w_0_170_s_0_540 = 2.87e-11  mcm2l1f_cf_w_0_170_s_0_540 = 2.03e-11
+ mcm2l1f_ca_w_0_170_s_0_720 = 9.12e-05  mcm2l1f_cc_w_0_170_s_0_720 = 1.96e-11  mcm2l1f_cf_w_0_170_s_0_720 = 2.53e-11
+ mcm2l1f_ca_w_0_170_s_1_080 = 9.12e-05  mcm2l1f_cc_w_0_170_s_1_080 = 9.80e-12  mcm2l1f_cf_w_0_170_s_1_080 = 3.22e-11
+ mcm2l1f_ca_w_0_170_s_1_980 = 9.12e-05  mcm2l1f_cc_w_0_170_s_1_980 = 1.89e-12  mcm2l1f_cf_w_0_170_s_1_980 = 3.91e-11
+ mcm2l1f_ca_w_0_170_s_4_500 = 9.12e-05  mcm2l1f_cc_w_0_170_s_4_500 = 5.00e-14  mcm2l1f_cf_w_0_170_s_4_500 = 4.09e-11
+ mcm2l1f_ca_w_1_360_s_0_180 = 9.12e-05  mcm2l1f_cc_w_1_360_s_0_180 = 9.40e-11  mcm2l1f_cf_w_1_360_s_0_180 = 6.90e-12
+ mcm2l1f_ca_w_1_360_s_0_225 = 9.12e-05  mcm2l1f_cc_w_1_360_s_0_225 = 7.63e-11  mcm2l1f_cf_w_1_360_s_0_225 = 8.80e-12
+ mcm2l1f_ca_w_1_360_s_0_270 = 9.12e-05  mcm2l1f_cc_w_1_360_s_0_270 = 6.43e-11  mcm2l1f_cf_w_1_360_s_0_270 = 1.06e-11
+ mcm2l1f_ca_w_1_360_s_0_360 = 9.12e-05  mcm2l1f_cc_w_1_360_s_0_360 = 4.88e-11  mcm2l1f_cf_w_1_360_s_0_360 = 1.42e-11
+ mcm2l1f_ca_w_1_360_s_0_450 = 9.12e-05  mcm2l1f_cc_w_1_360_s_0_450 = 3.86e-11  mcm2l1f_cf_w_1_360_s_0_450 = 1.74e-11
+ mcm2l1f_ca_w_1_360_s_0_540 = 9.12e-05  mcm2l1f_cc_w_1_360_s_0_540 = 3.14e-11  mcm2l1f_cf_w_1_360_s_0_540 = 2.04e-11
+ mcm2l1f_ca_w_1_360_s_0_720 = 9.12e-05  mcm2l1f_cc_w_1_360_s_0_720 = 2.15e-11  mcm2l1f_cf_w_1_360_s_0_720 = 2.56e-11
+ mcm2l1f_ca_w_1_360_s_1_080 = 9.12e-05  mcm2l1f_cc_w_1_360_s_1_080 = 1.08e-11  mcm2l1f_cf_w_1_360_s_1_080 = 3.30e-11
+ mcm2l1f_ca_w_1_360_s_1_980 = 9.12e-05  mcm2l1f_cc_w_1_360_s_1_980 = 2.20e-12  mcm2l1f_cf_w_1_360_s_1_980 = 4.05e-11
+ mcm2l1f_ca_w_1_360_s_4_500 = 9.12e-05  mcm2l1f_cc_w_1_360_s_4_500 = 0.00e+00  mcm2l1f_cf_w_1_360_s_4_500 = 4.26e-11
+ mcm2l1d_ca_w_0_170_s_0_180 = 1.12e-04  mcm2l1d_cc_w_0_170_s_0_180 = 8.44e-11  mcm2l1d_cf_w_0_170_s_0_180 = 8.45e-12
+ mcm2l1d_ca_w_0_170_s_0_225 = 1.12e-04  mcm2l1d_cc_w_0_170_s_0_225 = 6.78e-11  mcm2l1d_cf_w_0_170_s_0_225 = 1.07e-11
+ mcm2l1d_ca_w_0_170_s_0_270 = 1.12e-04  mcm2l1d_cc_w_0_170_s_0_270 = 5.63e-11  mcm2l1d_cf_w_0_170_s_0_270 = 1.29e-11
+ mcm2l1d_ca_w_0_170_s_0_360 = 1.12e-04  mcm2l1d_cc_w_0_170_s_0_360 = 4.17e-11  mcm2l1d_cf_w_0_170_s_0_360 = 1.71e-11
+ mcm2l1d_ca_w_0_170_s_0_450 = 1.12e-04  mcm2l1d_cc_w_0_170_s_0_450 = 3.23e-11  mcm2l1d_cf_w_0_170_s_0_450 = 2.08e-11
+ mcm2l1d_ca_w_0_170_s_0_540 = 1.12e-04  mcm2l1d_cc_w_0_170_s_0_540 = 2.56e-11  mcm2l1d_cf_w_0_170_s_0_540 = 2.41e-11
+ mcm2l1d_ca_w_0_170_s_0_720 = 1.12e-04  mcm2l1d_cc_w_0_170_s_0_720 = 1.66e-11  mcm2l1d_cf_w_0_170_s_0_720 = 2.95e-11
+ mcm2l1d_ca_w_0_170_s_1_080 = 1.12e-04  mcm2l1d_cc_w_0_170_s_1_080 = 7.51e-12  mcm2l1d_cf_w_0_170_s_1_080 = 3.65e-11
+ mcm2l1d_ca_w_0_170_s_1_980 = 1.12e-04  mcm2l1d_cc_w_0_170_s_1_980 = 1.13e-12  mcm2l1d_cf_w_0_170_s_1_980 = 4.24e-11
+ mcm2l1d_ca_w_0_170_s_4_500 = 1.12e-04  mcm2l1d_cc_w_0_170_s_4_500 = 4.50e-14  mcm2l1d_cf_w_0_170_s_4_500 = 4.35e-11
+ mcm2l1d_ca_w_1_360_s_0_180 = 1.12e-04  mcm2l1d_cc_w_1_360_s_0_180 = 9.01e-11  mcm2l1d_cf_w_1_360_s_0_180 = 8.42e-12
+ mcm2l1d_ca_w_1_360_s_0_225 = 1.12e-04  mcm2l1d_cc_w_1_360_s_0_225 = 7.23e-11  mcm2l1d_cf_w_1_360_s_0_225 = 1.07e-11
+ mcm2l1d_ca_w_1_360_s_0_270 = 1.12e-04  mcm2l1d_cc_w_1_360_s_0_270 = 6.03e-11  mcm2l1d_cf_w_1_360_s_0_270 = 1.29e-11
+ mcm2l1d_ca_w_1_360_s_0_360 = 1.12e-04  mcm2l1d_cc_w_1_360_s_0_360 = 4.48e-11  mcm2l1d_cf_w_1_360_s_0_360 = 1.71e-11
+ mcm2l1d_ca_w_1_360_s_0_450 = 1.12e-04  mcm2l1d_cc_w_1_360_s_0_450 = 3.47e-11  mcm2l1d_cf_w_1_360_s_0_450 = 2.09e-11
+ mcm2l1d_ca_w_1_360_s_0_540 = 1.12e-04  mcm2l1d_cc_w_1_360_s_0_540 = 2.75e-11  mcm2l1d_cf_w_1_360_s_0_540 = 2.43e-11
+ mcm2l1d_ca_w_1_360_s_0_720 = 1.12e-04  mcm2l1d_cc_w_1_360_s_0_720 = 1.80e-11  mcm2l1d_cf_w_1_360_s_0_720 = 2.99e-11
+ mcm2l1d_ca_w_1_360_s_1_080 = 1.12e-04  mcm2l1d_cc_w_1_360_s_1_080 = 8.28e-12  mcm2l1d_cf_w_1_360_s_1_080 = 3.73e-11
+ mcm2l1d_ca_w_1_360_s_1_980 = 1.12e-04  mcm2l1d_cc_w_1_360_s_1_980 = 1.28e-12  mcm2l1d_cf_w_1_360_s_1_980 = 4.37e-11
+ mcm2l1d_ca_w_1_360_s_4_500 = 1.12e-04  mcm2l1d_cc_w_1_360_s_4_500 = 5.00e-14  mcm2l1d_cf_w_1_360_s_4_500 = 4.49e-11
+ mcm2l1p1_ca_w_0_170_s_0_180 = 1.86e-04  mcm2l1p1_cc_w_0_170_s_0_180 = 7.79e-11  mcm2l1p1_cf_w_0_170_s_0_180 = 1.37e-11
+ mcm2l1p1_ca_w_0_170_s_0_225 = 1.86e-04  mcm2l1p1_cc_w_0_170_s_0_225 = 6.08e-11  mcm2l1p1_cf_w_0_170_s_0_225 = 1.73e-11
+ mcm2l1p1_ca_w_0_170_s_0_270 = 1.86e-04  mcm2l1p1_cc_w_0_170_s_0_270 = 4.94e-11  mcm2l1p1_cf_w_0_170_s_0_270 = 2.06e-11
+ mcm2l1p1_ca_w_0_170_s_0_360 = 1.86e-04  mcm2l1p1_cc_w_0_170_s_0_360 = 3.46e-11  mcm2l1p1_cf_w_0_170_s_0_360 = 2.66e-11
+ mcm2l1p1_ca_w_0_170_s_0_450 = 1.86e-04  mcm2l1p1_cc_w_0_170_s_0_450 = 2.54e-11  mcm2l1p1_cf_w_0_170_s_0_450 = 3.15e-11
+ mcm2l1p1_ca_w_0_170_s_0_540 = 1.86e-04  mcm2l1p1_cc_w_0_170_s_0_540 = 1.90e-11  mcm2l1p1_cf_w_0_170_s_0_540 = 3.57e-11
+ mcm2l1p1_ca_w_0_170_s_0_720 = 1.86e-04  mcm2l1p1_cc_w_0_170_s_0_720 = 1.10e-11  mcm2l1p1_cf_w_0_170_s_0_720 = 4.17e-11
+ mcm2l1p1_ca_w_0_170_s_1_080 = 1.86e-04  mcm2l1p1_cc_w_0_170_s_1_080 = 3.99e-12  mcm2l1p1_cf_w_0_170_s_1_080 = 4.79e-11
+ mcm2l1p1_ca_w_0_170_s_1_980 = 1.86e-04  mcm2l1p1_cc_w_0_170_s_1_980 = 3.90e-13  mcm2l1p1_cf_w_0_170_s_1_980 = 5.13e-11
+ mcm2l1p1_ca_w_0_170_s_4_500 = 1.86e-04  mcm2l1p1_cc_w_0_170_s_4_500 = 3.50e-14  mcm2l1p1_cf_w_0_170_s_4_500 = 5.17e-11
+ mcm2l1p1_ca_w_1_360_s_0_180 = 1.86e-04  mcm2l1p1_cc_w_1_360_s_0_180 = 8.20e-11  mcm2l1p1_cf_w_1_360_s_0_180 = 1.37e-11
+ mcm2l1p1_ca_w_1_360_s_0_225 = 1.86e-04  mcm2l1p1_cc_w_1_360_s_0_225 = 6.42e-11  mcm2l1p1_cf_w_1_360_s_0_225 = 1.72e-11
+ mcm2l1p1_ca_w_1_360_s_0_270 = 1.86e-04  mcm2l1p1_cc_w_1_360_s_0_270 = 5.24e-11  mcm2l1p1_cf_w_1_360_s_0_270 = 2.05e-11
+ mcm2l1p1_ca_w_1_360_s_0_360 = 1.86e-04  mcm2l1p1_cc_w_1_360_s_0_360 = 3.70e-11  mcm2l1p1_cf_w_1_360_s_0_360 = 2.65e-11
+ mcm2l1p1_ca_w_1_360_s_0_450 = 1.86e-04  mcm2l1p1_cc_w_1_360_s_0_450 = 2.73e-11  mcm2l1p1_cf_w_1_360_s_0_450 = 3.16e-11
+ mcm2l1p1_ca_w_1_360_s_0_540 = 1.86e-04  mcm2l1p1_cc_w_1_360_s_0_540 = 2.06e-11  mcm2l1p1_cf_w_1_360_s_0_540 = 3.58e-11
+ mcm2l1p1_ca_w_1_360_s_0_720 = 1.86e-04  mcm2l1p1_cc_w_1_360_s_0_720 = 1.21e-11  mcm2l1p1_cf_w_1_360_s_0_720 = 4.21e-11
+ mcm2l1p1_ca_w_1_360_s_1_080 = 1.86e-04  mcm2l1p1_cc_w_1_360_s_1_080 = 4.45e-12  mcm2l1p1_cf_w_1_360_s_1_080 = 4.87e-11
+ mcm2l1p1_ca_w_1_360_s_1_980 = 1.86e-04  mcm2l1p1_cc_w_1_360_s_1_980 = 4.25e-13  mcm2l1p1_cf_w_1_360_s_1_980 = 5.26e-11
+ mcm2l1p1_ca_w_1_360_s_4_500 = 1.86e-04  mcm2l1p1_cc_w_1_360_s_4_500 = 1.00e-14  mcm2l1p1_cf_w_1_360_s_4_500 = 5.29e-11
+ mcm3l1f_ca_w_0_170_s_0_180 = 6.92e-05  mcm3l1f_cc_w_0_170_s_0_180 = 9.00e-11  mcm3l1f_cf_w_0_170_s_0_180 = 5.30e-12
+ mcm3l1f_ca_w_0_170_s_0_225 = 6.92e-05  mcm3l1f_cc_w_0_170_s_0_225 = 7.36e-11  mcm3l1f_cf_w_0_170_s_0_225 = 6.76e-12
+ mcm3l1f_ca_w_0_170_s_0_270 = 6.92e-05  mcm3l1f_cc_w_0_170_s_0_270 = 6.28e-11  mcm3l1f_cf_w_0_170_s_0_270 = 8.19e-12
+ mcm3l1f_ca_w_0_170_s_0_360 = 6.92e-05  mcm3l1f_cc_w_0_170_s_0_360 = 4.85e-11  mcm3l1f_cf_w_0_170_s_0_360 = 1.11e-11
+ mcm3l1f_ca_w_0_170_s_0_450 = 6.92e-05  mcm3l1f_cc_w_0_170_s_0_450 = 3.96e-11  mcm3l1f_cf_w_0_170_s_0_450 = 1.35e-11
+ mcm3l1f_ca_w_0_170_s_0_540 = 6.92e-05  mcm3l1f_cc_w_0_170_s_0_540 = 3.30e-11  mcm3l1f_cf_w_0_170_s_0_540 = 1.60e-11
+ mcm3l1f_ca_w_0_170_s_0_720 = 6.92e-05  mcm3l1f_cc_w_0_170_s_0_720 = 2.40e-11  mcm3l1f_cf_w_0_170_s_0_720 = 2.03e-11
+ mcm3l1f_ca_w_0_170_s_1_080 = 6.92e-05  mcm3l1f_cc_w_0_170_s_1_080 = 1.37e-11  mcm3l1f_cf_w_0_170_s_1_080 = 2.67e-11
+ mcm3l1f_ca_w_0_170_s_1_980 = 6.92e-05  mcm3l1f_cc_w_0_170_s_1_980 = 3.89e-12  mcm3l1f_cf_w_0_170_s_1_980 = 3.47e-11
+ mcm3l1f_ca_w_0_170_s_4_500 = 6.92e-05  mcm3l1f_cc_w_0_170_s_4_500 = 1.75e-13  mcm3l1f_cf_w_0_170_s_4_500 = 3.82e-11
+ mcm3l1f_ca_w_1_360_s_0_180 = 6.92e-05  mcm3l1f_cc_w_1_360_s_0_180 = 1.01e-10  mcm3l1f_cf_w_1_360_s_0_180 = 5.28e-12
+ mcm3l1f_ca_w_1_360_s_0_225 = 6.92e-05  mcm3l1f_cc_w_1_360_s_0_225 = 8.31e-11  mcm3l1f_cf_w_1_360_s_0_225 = 6.75e-12
+ mcm3l1f_ca_w_1_360_s_0_270 = 6.92e-05  mcm3l1f_cc_w_1_360_s_0_270 = 7.12e-11  mcm3l1f_cf_w_1_360_s_0_270 = 8.19e-12
+ mcm3l1f_ca_w_1_360_s_0_360 = 6.92e-05  mcm3l1f_cc_w_1_360_s_0_360 = 5.56e-11  mcm3l1f_cf_w_1_360_s_0_360 = 1.10e-11
+ mcm3l1f_ca_w_1_360_s_0_450 = 6.92e-05  mcm3l1f_cc_w_1_360_s_0_450 = 4.54e-11  mcm3l1f_cf_w_1_360_s_0_450 = 1.36e-11
+ mcm3l1f_ca_w_1_360_s_0_540 = 6.92e-05  mcm3l1f_cc_w_1_360_s_0_540 = 3.80e-11  mcm3l1f_cf_w_1_360_s_0_540 = 1.61e-11
+ mcm3l1f_ca_w_1_360_s_0_720 = 6.92e-05  mcm3l1f_cc_w_1_360_s_0_720 = 2.78e-11  mcm3l1f_cf_w_1_360_s_0_720 = 2.05e-11
+ mcm3l1f_ca_w_1_360_s_1_080 = 6.92e-05  mcm3l1f_cc_w_1_360_s_1_080 = 1.62e-11  mcm3l1f_cf_w_1_360_s_1_080 = 2.74e-11
+ mcm3l1f_ca_w_1_360_s_1_980 = 6.92e-05  mcm3l1f_cc_w_1_360_s_1_980 = 4.77e-12  mcm3l1f_cf_w_1_360_s_1_980 = 3.66e-11
+ mcm3l1f_ca_w_1_360_s_4_500 = 6.92e-05  mcm3l1f_cc_w_1_360_s_4_500 = 2.25e-13  mcm3l1f_cf_w_1_360_s_4_500 = 4.09e-11
+ mcm3l1d_ca_w_0_170_s_0_180 = 8.97e-05  mcm3l1d_cc_w_0_170_s_0_180 = 8.75e-11  mcm3l1d_cf_w_0_170_s_0_180 = 6.82e-12
+ mcm3l1d_ca_w_0_170_s_0_225 = 8.97e-05  mcm3l1d_cc_w_0_170_s_0_225 = 7.10e-11  mcm3l1d_cf_w_0_170_s_0_225 = 8.68e-12
+ mcm3l1d_ca_w_0_170_s_0_270 = 8.97e-05  mcm3l1d_cc_w_0_170_s_0_270 = 6.00e-11  mcm3l1d_cf_w_0_170_s_0_270 = 1.05e-11
+ mcm3l1d_ca_w_0_170_s_0_360 = 8.97e-05  mcm3l1d_cc_w_0_170_s_0_360 = 4.55e-11  mcm3l1d_cf_w_0_170_s_0_360 = 1.40e-11
+ mcm3l1d_ca_w_0_170_s_0_450 = 8.97e-05  mcm3l1d_cc_w_0_170_s_0_450 = 3.64e-11  mcm3l1d_cf_w_0_170_s_0_450 = 1.71e-11
+ mcm3l1d_ca_w_0_170_s_0_540 = 8.97e-05  mcm3l1d_cc_w_0_170_s_0_540 = 2.97e-11  mcm3l1d_cf_w_0_170_s_0_540 = 2.01e-11
+ mcm3l1d_ca_w_0_170_s_0_720 = 8.97e-05  mcm3l1d_cc_w_0_170_s_0_720 = 2.08e-11  mcm3l1d_cf_w_0_170_s_0_720 = 2.49e-11
+ mcm3l1d_ca_w_0_170_s_1_080 = 8.97e-05  mcm3l1d_cc_w_0_170_s_1_080 = 1.10e-11  mcm3l1d_cf_w_0_170_s_1_080 = 3.18e-11
+ mcm3l1d_ca_w_0_170_s_1_980 = 8.97e-05  mcm3l1d_cc_w_0_170_s_1_980 = 2.64e-12  mcm3l1d_cf_w_0_170_s_1_980 = 3.90e-11
+ mcm3l1d_ca_w_0_170_s_4_500 = 8.97e-05  mcm3l1d_cc_w_0_170_s_4_500 = 9.50e-14  mcm3l1d_cf_w_0_170_s_4_500 = 4.15e-11
+ mcm3l1d_ca_w_1_360_s_0_180 = 8.97e-05  mcm3l1d_cc_w_1_360_s_0_180 = 9.66e-11  mcm3l1d_cf_w_1_360_s_0_180 = 6.80e-12
+ mcm3l1d_ca_w_1_360_s_0_225 = 8.97e-05  mcm3l1d_cc_w_1_360_s_0_225 = 7.89e-11  mcm3l1d_cf_w_1_360_s_0_225 = 8.67e-12
+ mcm3l1d_ca_w_1_360_s_0_270 = 8.97e-05  mcm3l1d_cc_w_1_360_s_0_270 = 6.71e-11  mcm3l1d_cf_w_1_360_s_0_270 = 1.05e-11
+ mcm3l1d_ca_w_1_360_s_0_360 = 8.97e-05  mcm3l1d_cc_w_1_360_s_0_360 = 5.15e-11  mcm3l1d_cf_w_1_360_s_0_360 = 1.39e-11
+ mcm3l1d_ca_w_1_360_s_0_450 = 8.97e-05  mcm3l1d_cc_w_1_360_s_0_450 = 4.13e-11  mcm3l1d_cf_w_1_360_s_0_450 = 1.72e-11
+ mcm3l1d_ca_w_1_360_s_0_540 = 8.97e-05  mcm3l1d_cc_w_1_360_s_0_540 = 3.40e-11  mcm3l1d_cf_w_1_360_s_0_540 = 2.01e-11
+ mcm3l1d_ca_w_1_360_s_0_720 = 8.97e-05  mcm3l1d_cc_w_1_360_s_0_720 = 2.41e-11  mcm3l1d_cf_w_1_360_s_0_720 = 2.52e-11
+ mcm3l1d_ca_w_1_360_s_1_080 = 8.97e-05  mcm3l1d_cc_w_1_360_s_1_080 = 1.31e-11  mcm3l1d_cf_w_1_360_s_1_080 = 3.27e-11
+ mcm3l1d_ca_w_1_360_s_1_980 = 8.97e-05  mcm3l1d_cc_w_1_360_s_1_980 = 3.28e-12  mcm3l1d_cf_w_1_360_s_1_980 = 4.11e-11
+ mcm3l1d_ca_w_1_360_s_4_500 = 8.97e-05  mcm3l1d_cc_w_1_360_s_4_500 = 1.60e-13  mcm3l1d_cf_w_1_360_s_4_500 = 4.41e-11
+ mcm3l1p1_ca_w_0_170_s_0_180 = 1.64e-04  mcm3l1p1_cc_w_0_170_s_0_180 = 8.10e-11  mcm3l1p1_cf_w_0_170_s_0_180 = 1.21e-11
+ mcm3l1p1_ca_w_0_170_s_0_225 = 1.64e-04  mcm3l1p1_cc_w_0_170_s_0_225 = 6.41e-11  mcm3l1p1_cf_w_0_170_s_0_225 = 1.53e-11
+ mcm3l1p1_ca_w_0_170_s_0_270 = 1.64e-04  mcm3l1p1_cc_w_0_170_s_0_270 = 5.29e-11  mcm3l1p1_cf_w_0_170_s_0_270 = 1.82e-11
+ mcm3l1p1_ca_w_0_170_s_0_360 = 1.64e-04  mcm3l1p1_cc_w_0_170_s_0_360 = 3.83e-11  mcm3l1p1_cf_w_0_170_s_0_360 = 2.38e-11
+ mcm3l1p1_ca_w_0_170_s_0_450 = 1.64e-04  mcm3l1p1_cc_w_0_170_s_0_450 = 2.93e-11  mcm3l1p1_cf_w_0_170_s_0_450 = 2.82e-11
+ mcm3l1p1_ca_w_0_170_s_0_540 = 1.64e-04  mcm3l1p1_cc_w_0_170_s_0_540 = 2.27e-11  mcm3l1p1_cf_w_0_170_s_0_540 = 3.22e-11
+ mcm3l1p1_ca_w_0_170_s_0_720 = 1.64e-04  mcm3l1p1_cc_w_0_170_s_0_720 = 1.45e-11  mcm3l1p1_cf_w_0_170_s_0_720 = 3.81e-11
+ mcm3l1p1_ca_w_0_170_s_1_080 = 1.64e-04  mcm3l1p1_cc_w_0_170_s_1_080 = 6.50e-12  mcm3l1p1_cf_w_0_170_s_1_080 = 4.48e-11
+ mcm3l1p1_ca_w_0_170_s_1_980 = 1.64e-04  mcm3l1p1_cc_w_0_170_s_1_980 = 1.18e-12  mcm3l1p1_cf_w_0_170_s_1_980 = 4.98e-11
+ mcm3l1p1_ca_w_0_170_s_4_500 = 1.64e-04  mcm3l1p1_cc_w_0_170_s_4_500 = 4.00e-14  mcm3l1p1_cf_w_0_170_s_4_500 = 5.09e-11
+ mcm3l1p1_ca_w_1_360_s_0_180 = 1.64e-04  mcm3l1p1_cc_w_1_360_s_0_180 = 8.87e-11  mcm3l1p1_cf_w_1_360_s_0_180 = 1.21e-11
+ mcm3l1p1_ca_w_1_360_s_0_225 = 1.64e-04  mcm3l1p1_cc_w_1_360_s_0_225 = 7.09e-11  mcm3l1p1_cf_w_1_360_s_0_225 = 1.52e-11
+ mcm3l1p1_ca_w_1_360_s_0_270 = 1.64e-04  mcm3l1p1_cc_w_1_360_s_0_270 = 5.91e-11  mcm3l1p1_cf_w_1_360_s_0_270 = 1.82e-11
+ mcm3l1p1_ca_w_1_360_s_0_360 = 1.64e-04  mcm3l1p1_cc_w_1_360_s_0_360 = 4.37e-11  mcm3l1p1_cf_w_1_360_s_0_360 = 2.36e-11
+ mcm3l1p1_ca_w_1_360_s_0_450 = 1.64e-04  mcm3l1p1_cc_w_1_360_s_0_450 = 3.37e-11  mcm3l1p1_cf_w_1_360_s_0_450 = 2.83e-11
+ mcm3l1p1_ca_w_1_360_s_0_540 = 1.64e-04  mcm3l1p1_cc_w_1_360_s_0_540 = 2.67e-11  mcm3l1p1_cf_w_1_360_s_0_540 = 3.23e-11
+ mcm3l1p1_ca_w_1_360_s_0_720 = 1.64e-04  mcm3l1p1_cc_w_1_360_s_0_720 = 1.76e-11  mcm3l1p1_cf_w_1_360_s_0_720 = 3.86e-11
+ mcm3l1p1_ca_w_1_360_s_1_080 = 1.64e-04  mcm3l1p1_cc_w_1_360_s_1_080 = 8.40e-12  mcm3l1p1_cf_w_1_360_s_1_080 = 4.62e-11
+ mcm3l1p1_ca_w_1_360_s_1_980 = 1.64e-04  mcm3l1p1_cc_w_1_360_s_1_980 = 1.62e-12  mcm3l1p1_cf_w_1_360_s_1_980 = 5.25e-11
+ mcm3l1p1_ca_w_1_360_s_4_500 = 1.64e-04  mcm3l1p1_cc_w_1_360_s_4_500 = 3.50e-14  mcm3l1p1_cf_w_1_360_s_4_500 = 5.40e-11
+ mcm4l1f_ca_w_0_170_s_0_180 = 5.85e-05  mcm4l1f_cc_w_0_170_s_0_180 = 9.15e-11  mcm4l1f_cf_w_0_170_s_0_180 = 4.49e-12
+ mcm4l1f_ca_w_0_170_s_0_225 = 5.85e-05  mcm4l1f_cc_w_0_170_s_0_225 = 7.52e-11  mcm4l1f_cf_w_0_170_s_0_225 = 5.74e-12
+ mcm4l1f_ca_w_0_170_s_0_270 = 5.85e-05  mcm4l1f_cc_w_0_170_s_0_270 = 6.48e-11  mcm4l1f_cf_w_0_170_s_0_270 = 6.96e-12
+ mcm4l1f_ca_w_0_170_s_0_360 = 5.85e-05  mcm4l1f_cc_w_0_170_s_0_360 = 5.08e-11  mcm4l1f_cf_w_0_170_s_0_360 = 9.47e-12
+ mcm4l1f_ca_w_0_170_s_0_450 = 5.85e-05  mcm4l1f_cc_w_0_170_s_0_450 = 4.21e-11  mcm4l1f_cf_w_0_170_s_0_450 = 1.16e-11
+ mcm4l1f_ca_w_0_170_s_0_540 = 5.85e-05  mcm4l1f_cc_w_0_170_s_0_540 = 3.56e-11  mcm4l1f_cf_w_0_170_s_0_540 = 1.38e-11
+ mcm4l1f_ca_w_0_170_s_0_720 = 5.85e-05  mcm4l1f_cc_w_0_170_s_0_720 = 2.68e-11  mcm4l1f_cf_w_0_170_s_0_720 = 1.76e-11
+ mcm4l1f_ca_w_0_170_s_1_080 = 5.85e-05  mcm4l1f_cc_w_0_170_s_1_080 = 1.65e-11  mcm4l1f_cf_w_0_170_s_1_080 = 2.36e-11
+ mcm4l1f_ca_w_0_170_s_1_980 = 5.85e-05  mcm4l1f_cc_w_0_170_s_1_980 = 5.98e-12  mcm4l1f_cf_w_0_170_s_1_980 = 3.18e-11
+ mcm4l1f_ca_w_0_170_s_4_500 = 5.85e-05  mcm4l1f_cc_w_0_170_s_4_500 = 5.45e-13  mcm4l1f_cf_w_0_170_s_4_500 = 3.68e-11
+ mcm4l1f_ca_w_1_360_s_0_180 = 5.85e-05  mcm4l1f_cc_w_1_360_s_0_180 = 1.06e-10  mcm4l1f_cf_w_1_360_s_0_180 = 4.49e-12
+ mcm4l1f_ca_w_1_360_s_0_225 = 5.85e-05  mcm4l1f_cc_w_1_360_s_0_225 = 8.82e-11  mcm4l1f_cf_w_1_360_s_0_225 = 5.74e-12
+ mcm4l1f_ca_w_1_360_s_0_270 = 5.85e-05  mcm4l1f_cc_w_1_360_s_0_270 = 7.63e-11  mcm4l1f_cf_w_1_360_s_0_270 = 6.97e-12
+ mcm4l1f_ca_w_1_360_s_0_360 = 5.85e-05  mcm4l1f_cc_w_1_360_s_0_360 = 6.08e-11  mcm4l1f_cf_w_1_360_s_0_360 = 9.34e-12
+ mcm4l1f_ca_w_1_360_s_0_450 = 5.85e-05  mcm4l1f_cc_w_1_360_s_0_450 = 5.05e-11  mcm4l1f_cf_w_1_360_s_0_450 = 1.16e-11
+ mcm4l1f_ca_w_1_360_s_0_540 = 5.85e-05  mcm4l1f_cc_w_1_360_s_0_540 = 4.32e-11  mcm4l1f_cf_w_1_360_s_0_540 = 1.38e-11
+ mcm4l1f_ca_w_1_360_s_0_720 = 5.85e-05  mcm4l1f_cc_w_1_360_s_0_720 = 3.30e-11  mcm4l1f_cf_w_1_360_s_0_720 = 1.77e-11
+ mcm4l1f_ca_w_1_360_s_1_080 = 5.85e-05  mcm4l1f_cc_w_1_360_s_1_080 = 2.10e-11  mcm4l1f_cf_w_1_360_s_1_080 = 2.42e-11
+ mcm4l1f_ca_w_1_360_s_1_980 = 5.85e-05  mcm4l1f_cc_w_1_360_s_1_980 = 8.12e-12  mcm4l1f_cf_w_1_360_s_1_980 = 3.38e-11
+ mcm4l1f_ca_w_1_360_s_4_500 = 5.85e-05  mcm4l1f_cc_w_1_360_s_4_500 = 7.90e-13  mcm4l1f_cf_w_1_360_s_4_500 = 4.06e-11
+ mcm4l1d_ca_w_0_170_s_0_180 = 7.90e-05  mcm4l1d_cc_w_0_170_s_0_180 = 8.91e-11  mcm4l1d_cf_w_0_170_s_0_180 = 6.02e-12
+ mcm4l1d_ca_w_0_170_s_0_225 = 7.90e-05  mcm4l1d_cc_w_0_170_s_0_225 = 7.25e-11  mcm4l1d_cf_w_0_170_s_0_225 = 7.66e-12
+ mcm4l1d_ca_w_0_170_s_0_270 = 7.90e-05  mcm4l1d_cc_w_0_170_s_0_270 = 6.19e-11  mcm4l1d_cf_w_0_170_s_0_270 = 9.26e-12
+ mcm4l1d_ca_w_0_170_s_0_360 = 7.90e-05  mcm4l1d_cc_w_0_170_s_0_360 = 4.77e-11  mcm4l1d_cf_w_0_170_s_0_360 = 1.25e-11
+ mcm4l1d_ca_w_0_170_s_0_450 = 7.90e-05  mcm4l1d_cc_w_0_170_s_0_450 = 3.88e-11  mcm4l1d_cf_w_0_170_s_0_450 = 1.52e-11
+ mcm4l1d_ca_w_0_170_s_0_540 = 7.90e-05  mcm4l1d_cc_w_0_170_s_0_540 = 3.22e-11  mcm4l1d_cf_w_0_170_s_0_540 = 1.80e-11
+ mcm4l1d_ca_w_0_170_s_0_720 = 7.90e-05  mcm4l1d_cc_w_0_170_s_0_720 = 2.34e-11  mcm4l1d_cf_w_0_170_s_0_720 = 2.25e-11
+ mcm4l1d_ca_w_0_170_s_1_080 = 7.90e-05  mcm4l1d_cc_w_0_170_s_1_080 = 1.35e-11  mcm4l1d_cf_w_0_170_s_1_080 = 2.91e-11
+ mcm4l1d_ca_w_0_170_s_1_980 = 7.90e-05  mcm4l1d_cc_w_0_170_s_1_980 = 4.27e-12  mcm4l1d_cf_w_0_170_s_1_980 = 3.69e-11
+ mcm4l1d_ca_w_0_170_s_4_500 = 7.90e-05  mcm4l1d_cc_w_0_170_s_4_500 = 3.25e-13  mcm4l1d_cf_w_0_170_s_4_500 = 4.06e-11
+ mcm4l1d_ca_w_1_360_s_0_180 = 7.90e-05  mcm4l1d_cc_w_1_360_s_0_180 = 1.02e-10  mcm4l1d_cf_w_1_360_s_0_180 = 6.01e-12
+ mcm4l1d_ca_w_1_360_s_0_225 = 7.90e-05  mcm4l1d_cc_w_1_360_s_0_225 = 8.40e-11  mcm4l1d_cf_w_1_360_s_0_225 = 7.66e-12
+ mcm4l1d_ca_w_1_360_s_0_270 = 7.90e-05  mcm4l1d_cc_w_1_360_s_0_270 = 7.22e-11  mcm4l1d_cf_w_1_360_s_0_270 = 9.26e-12
+ mcm4l1d_ca_w_1_360_s_0_360 = 7.90e-05  mcm4l1d_cc_w_1_360_s_0_360 = 5.67e-11  mcm4l1d_cf_w_1_360_s_0_360 = 1.23e-11
+ mcm4l1d_ca_w_1_360_s_0_450 = 7.90e-05  mcm4l1d_cc_w_1_360_s_0_450 = 4.65e-11  mcm4l1d_cf_w_1_360_s_0_450 = 1.53e-11
+ mcm4l1d_ca_w_1_360_s_0_540 = 7.90e-05  mcm4l1d_cc_w_1_360_s_0_540 = 3.93e-11  mcm4l1d_cf_w_1_360_s_0_540 = 1.79e-11
+ mcm4l1d_ca_w_1_360_s_0_720 = 7.90e-05  mcm4l1d_cc_w_1_360_s_0_720 = 2.92e-11  mcm4l1d_cf_w_1_360_s_0_720 = 2.27e-11
+ mcm4l1d_ca_w_1_360_s_1_080 = 7.90e-05  mcm4l1d_cc_w_1_360_s_1_080 = 1.77e-11  mcm4l1d_cf_w_1_360_s_1_080 = 2.99e-11
+ mcm4l1d_ca_w_1_360_s_1_980 = 7.90e-05  mcm4l1d_cc_w_1_360_s_1_980 = 6.14e-12  mcm4l1d_cf_w_1_360_s_1_980 = 3.93e-11
+ mcm4l1d_ca_w_1_360_s_4_500 = 7.90e-05  mcm4l1d_cc_w_1_360_s_4_500 = 4.85e-13  mcm4l1d_cf_w_1_360_s_4_500 = 4.47e-11
+ mcm4l1p1_ca_w_0_170_s_0_180 = 1.53e-04  mcm4l1p1_cc_w_0_170_s_0_180 = 8.24e-11  mcm4l1p1_cf_w_0_170_s_0_180 = 1.13e-11
+ mcm4l1p1_ca_w_0_170_s_0_225 = 1.53e-04  mcm4l1p1_cc_w_0_170_s_0_225 = 6.57e-11  mcm4l1p1_cf_w_0_170_s_0_225 = 1.43e-11
+ mcm4l1p1_ca_w_0_170_s_0_270 = 1.53e-04  mcm4l1p1_cc_w_0_170_s_0_270 = 5.49e-11  mcm4l1p1_cf_w_0_170_s_0_270 = 1.70e-11
+ mcm4l1p1_ca_w_0_170_s_0_360 = 1.53e-04  mcm4l1p1_cc_w_0_170_s_0_360 = 4.03e-11  mcm4l1p1_cf_w_0_170_s_0_360 = 2.24e-11
+ mcm4l1p1_ca_w_0_170_s_0_450 = 1.53e-04  mcm4l1p1_cc_w_0_170_s_0_450 = 3.16e-11  mcm4l1p1_cf_w_0_170_s_0_450 = 2.65e-11
+ mcm4l1p1_ca_w_0_170_s_0_540 = 1.53e-04  mcm4l1p1_cc_w_0_170_s_0_540 = 2.49e-11  mcm4l1p1_cf_w_0_170_s_0_540 = 3.05e-11
+ mcm4l1p1_ca_w_0_170_s_0_720 = 1.53e-04  mcm4l1p1_cc_w_0_170_s_0_720 = 1.66e-11  mcm4l1p1_cf_w_0_170_s_0_720 = 3.63e-11
+ mcm4l1p1_ca_w_0_170_s_1_080 = 1.53e-04  mcm4l1p1_cc_w_0_170_s_1_080 = 8.37e-12  mcm4l1p1_cf_w_0_170_s_1_080 = 4.31e-11
+ mcm4l1p1_ca_w_0_170_s_1_980 = 1.53e-04  mcm4l1p1_cc_w_0_170_s_1_980 = 2.16e-12  mcm4l1p1_cf_w_0_170_s_1_980 = 4.89e-11
+ mcm4l1p1_ca_w_0_170_s_4_500 = 1.53e-04  mcm4l1p1_cc_w_0_170_s_4_500 = 1.50e-13  mcm4l1p1_cf_w_0_170_s_4_500 = 5.08e-11
+ mcm4l1p1_ca_w_1_360_s_0_180 = 1.53e-04  mcm4l1p1_cc_w_1_360_s_0_180 = 9.37e-11  mcm4l1p1_cf_w_1_360_s_0_180 = 1.15e-11
+ mcm4l1p1_ca_w_1_360_s_0_225 = 1.53e-04  mcm4l1p1_cc_w_1_360_s_0_225 = 7.62e-11  mcm4l1p1_cf_w_1_360_s_0_225 = 1.44e-11
+ mcm4l1p1_ca_w_1_360_s_0_270 = 1.53e-04  mcm4l1p1_cc_w_1_360_s_0_270 = 6.42e-11  mcm4l1p1_cf_w_1_360_s_0_270 = 1.72e-11
+ mcm4l1p1_ca_w_1_360_s_0_360 = 1.53e-04  mcm4l1p1_cc_w_1_360_s_0_360 = 4.88e-11  mcm4l1p1_cf_w_1_360_s_0_360 = 2.23e-11
+ mcm4l1p1_ca_w_1_360_s_0_450 = 1.53e-04  mcm4l1p1_cc_w_1_360_s_0_450 = 3.89e-11  mcm4l1p1_cf_w_1_360_s_0_450 = 2.67e-11
+ mcm4l1p1_ca_w_1_360_s_0_540 = 1.53e-04  mcm4l1p1_cc_w_1_360_s_0_540 = 3.18e-11  mcm4l1p1_cf_w_1_360_s_0_540 = 3.06e-11
+ mcm4l1p1_ca_w_1_360_s_0_720 = 1.53e-04  mcm4l1p1_cc_w_1_360_s_0_720 = 2.24e-11  mcm4l1p1_cf_w_1_360_s_0_720 = 3.68e-11
+ mcm4l1p1_ca_w_1_360_s_1_080 = 1.53e-04  mcm4l1p1_cc_w_1_360_s_1_080 = 1.24e-11  mcm4l1p1_cf_w_1_360_s_1_080 = 4.47e-11
+ mcm4l1p1_ca_w_1_360_s_1_980 = 1.53e-04  mcm4l1p1_cc_w_1_360_s_1_980 = 3.73e-12  mcm4l1p1_cf_w_1_360_s_1_980 = 5.25e-11
+ mcm4l1p1_ca_w_1_360_s_4_500 = 1.53e-04  mcm4l1p1_cc_w_1_360_s_4_500 = 2.90e-13  mcm4l1p1_cf_w_1_360_s_4_500 = 5.59e-11
+ mcm5l1f_ca_w_0_170_s_0_180 = 5.41e-05  mcm5l1f_cc_w_0_170_s_0_180 = 9.21e-11  mcm5l1f_cf_w_0_170_s_0_180 = 4.16e-12
+ mcm5l1f_ca_w_0_170_s_0_225 = 5.41e-05  mcm5l1f_cc_w_0_170_s_0_225 = 7.60e-11  mcm5l1f_cf_w_0_170_s_0_225 = 5.31e-12
+ mcm5l1f_ca_w_0_170_s_0_270 = 5.41e-05  mcm5l1f_cc_w_0_170_s_0_270 = 6.56e-11  mcm5l1f_cf_w_0_170_s_0_270 = 6.44e-12
+ mcm5l1f_ca_w_0_170_s_0_360 = 5.41e-05  mcm5l1f_cc_w_0_170_s_0_360 = 5.17e-11  mcm5l1f_cf_w_0_170_s_0_360 = 8.80e-12
+ mcm5l1f_ca_w_0_170_s_0_450 = 5.41e-05  mcm5l1f_cc_w_0_170_s_0_450 = 4.31e-11  mcm5l1f_cf_w_0_170_s_0_450 = 1.07e-11
+ mcm5l1f_ca_w_0_170_s_0_540 = 5.41e-05  mcm5l1f_cc_w_0_170_s_0_540 = 3.67e-11  mcm5l1f_cf_w_0_170_s_0_540 = 1.29e-11
+ mcm5l1f_ca_w_0_170_s_0_720 = 5.41e-05  mcm5l1f_cc_w_0_170_s_0_720 = 2.80e-11  mcm5l1f_cf_w_0_170_s_0_720 = 1.65e-11
+ mcm5l1f_ca_w_0_170_s_1_080 = 5.41e-05  mcm5l1f_cc_w_0_170_s_1_080 = 1.79e-11  mcm5l1f_cf_w_0_170_s_1_080 = 2.23e-11
+ mcm5l1f_ca_w_0_170_s_1_980 = 5.41e-05  mcm5l1f_cc_w_0_170_s_1_980 = 7.22e-12  mcm5l1f_cf_w_0_170_s_1_980 = 3.04e-11
+ mcm5l1f_ca_w_0_170_s_4_500 = 5.41e-05  mcm5l1f_cc_w_0_170_s_4_500 = 9.75e-13  mcm5l1f_cf_w_0_170_s_4_500 = 3.61e-11
+ mcm5l1f_ca_w_1_360_s_0_180 = 5.41e-05  mcm5l1f_cc_w_1_360_s_0_180 = 1.08e-10  mcm5l1f_cf_w_1_360_s_0_180 = 4.15e-12
+ mcm5l1f_ca_w_1_360_s_0_225 = 5.41e-05  mcm5l1f_cc_w_1_360_s_0_225 = 9.08e-11  mcm5l1f_cf_w_1_360_s_0_225 = 5.31e-12
+ mcm5l1f_ca_w_1_360_s_0_270 = 5.41e-05  mcm5l1f_cc_w_1_360_s_0_270 = 7.89e-11  mcm5l1f_cf_w_1_360_s_0_270 = 6.45e-12
+ mcm5l1f_ca_w_1_360_s_0_360 = 5.41e-05  mcm5l1f_cc_w_1_360_s_0_360 = 6.34e-11  mcm5l1f_cf_w_1_360_s_0_360 = 8.66e-12
+ mcm5l1f_ca_w_1_360_s_0_450 = 5.41e-05  mcm5l1f_cc_w_1_360_s_0_450 = 5.33e-11  mcm5l1f_cf_w_1_360_s_0_450 = 1.08e-11
+ mcm5l1f_ca_w_1_360_s_0_540 = 5.41e-05  mcm5l1f_cc_w_1_360_s_0_540 = 4.60e-11  mcm5l1f_cf_w_1_360_s_0_540 = 1.28e-11
+ mcm5l1f_ca_w_1_360_s_0_720 = 5.41e-05  mcm5l1f_cc_w_1_360_s_0_720 = 3.59e-11  mcm5l1f_cf_w_1_360_s_0_720 = 1.65e-11
+ mcm5l1f_ca_w_1_360_s_1_080 = 5.41e-05  mcm5l1f_cc_w_1_360_s_1_080 = 2.39e-11  mcm5l1f_cf_w_1_360_s_1_080 = 2.27e-11
+ mcm5l1f_ca_w_1_360_s_1_980 = 5.41e-05  mcm5l1f_cc_w_1_360_s_1_980 = 1.05e-11  mcm5l1f_cf_w_1_360_s_1_980 = 3.24e-11
+ mcm5l1f_ca_w_1_360_s_4_500 = 5.41e-05  mcm5l1f_cc_w_1_360_s_4_500 = 1.60e-12  mcm5l1f_cf_w_1_360_s_4_500 = 4.04e-11
+ mcm5l1d_ca_w_0_170_s_0_180 = 7.46e-05  mcm5l1d_cc_w_0_170_s_0_180 = 8.97e-11  mcm5l1d_cf_w_0_170_s_0_180 = 5.68e-12
+ mcm5l1d_ca_w_0_170_s_0_225 = 7.46e-05  mcm5l1d_cc_w_0_170_s_0_225 = 7.33e-11  mcm5l1d_cf_w_0_170_s_0_225 = 7.24e-12
+ mcm5l1d_ca_w_0_170_s_0_270 = 7.46e-05  mcm5l1d_cc_w_0_170_s_0_270 = 6.27e-11  mcm5l1d_cf_w_0_170_s_0_270 = 8.75e-12
+ mcm5l1d_ca_w_0_170_s_0_360 = 7.46e-05  mcm5l1d_cc_w_0_170_s_0_360 = 4.84e-11  mcm5l1d_cf_w_0_170_s_0_360 = 1.18e-11
+ mcm5l1d_ca_w_0_170_s_0_450 = 7.46e-05  mcm5l1d_cc_w_0_170_s_0_450 = 3.99e-11  mcm5l1d_cf_w_0_170_s_0_450 = 1.43e-11
+ mcm5l1d_ca_w_0_170_s_0_540 = 7.46e-05  mcm5l1d_cc_w_0_170_s_0_540 = 3.32e-11  mcm5l1d_cf_w_0_170_s_0_540 = 1.71e-11
+ mcm5l1d_ca_w_0_170_s_0_720 = 7.46e-05  mcm5l1d_cc_w_0_170_s_0_720 = 2.45e-11  mcm5l1d_cf_w_0_170_s_0_720 = 2.15e-11
+ mcm5l1d_ca_w_0_170_s_1_080 = 7.46e-05  mcm5l1d_cc_w_0_170_s_1_080 = 1.47e-11  mcm5l1d_cf_w_0_170_s_1_080 = 2.80e-11
+ mcm5l1d_ca_w_0_170_s_1_980 = 7.46e-05  mcm5l1d_cc_w_0_170_s_1_980 = 5.26e-12  mcm5l1d_cf_w_0_170_s_1_980 = 3.58e-11
+ mcm5l1d_ca_w_0_170_s_4_500 = 7.46e-05  mcm5l1d_cc_w_0_170_s_4_500 = 6.20e-13  mcm5l1d_cf_w_0_170_s_4_500 = 4.03e-11
+ mcm5l1d_ca_w_1_360_s_0_180 = 7.46e-05  mcm5l1d_cc_w_1_360_s_0_180 = 1.04e-10  mcm5l1d_cf_w_1_360_s_0_180 = 5.68e-12
+ mcm5l1d_ca_w_1_360_s_0_225 = 7.46e-05  mcm5l1d_cc_w_1_360_s_0_225 = 8.66e-11  mcm5l1d_cf_w_1_360_s_0_225 = 7.24e-12
+ mcm5l1d_ca_w_1_360_s_0_270 = 7.46e-05  mcm5l1d_cc_w_1_360_s_0_270 = 7.47e-11  mcm5l1d_cf_w_1_360_s_0_270 = 8.76e-12
+ mcm5l1d_ca_w_1_360_s_0_360 = 7.46e-05  mcm5l1d_cc_w_1_360_s_0_360 = 5.93e-11  mcm5l1d_cf_w_1_360_s_0_360 = 1.17e-11
+ mcm5l1d_ca_w_1_360_s_0_450 = 7.46e-05  mcm5l1d_cc_w_1_360_s_0_450 = 4.93e-11  mcm5l1d_cf_w_1_360_s_0_450 = 1.44e-11
+ mcm5l1d_ca_w_1_360_s_0_540 = 7.46e-05  mcm5l1d_cc_w_1_360_s_0_540 = 4.20e-11  mcm5l1d_cf_w_1_360_s_0_540 = 1.70e-11
+ mcm5l1d_ca_w_1_360_s_0_720 = 7.46e-05  mcm5l1d_cc_w_1_360_s_0_720 = 3.21e-11  mcm5l1d_cf_w_1_360_s_0_720 = 2.15e-11
+ mcm5l1d_ca_w_1_360_s_1_080 = 7.46e-05  mcm5l1d_cc_w_1_360_s_1_080 = 2.04e-11  mcm5l1d_cf_w_1_360_s_1_080 = 2.86e-11
+ mcm5l1d_ca_w_1_360_s_1_980 = 7.46e-05  mcm5l1d_cc_w_1_360_s_1_980 = 8.23e-12  mcm5l1d_cf_w_1_360_s_1_980 = 3.84e-11
+ mcm5l1d_ca_w_1_360_s_4_500 = 7.46e-05  mcm5l1d_cc_w_1_360_s_4_500 = 1.13e-12  mcm5l1d_cf_w_1_360_s_4_500 = 4.51e-11
+ mcm5l1p1_ca_w_0_170_s_0_180 = 1.49e-04  mcm5l1p1_cc_w_0_170_s_0_180 = 8.31e-11  mcm5l1p1_cf_w_0_170_s_0_180 = 1.10e-11
+ mcm5l1p1_ca_w_0_170_s_0_225 = 1.49e-04  mcm5l1p1_cc_w_0_170_s_0_225 = 6.64e-11  mcm5l1p1_cf_w_0_170_s_0_225 = 1.39e-11
+ mcm5l1p1_ca_w_0_170_s_0_270 = 1.49e-04  mcm5l1p1_cc_w_0_170_s_0_270 = 5.56e-11  mcm5l1p1_cf_w_0_170_s_0_270 = 1.65e-11
+ mcm5l1p1_ca_w_0_170_s_0_360 = 1.49e-04  mcm5l1p1_cc_w_0_170_s_0_360 = 4.11e-11  mcm5l1p1_cf_w_0_170_s_0_360 = 2.18e-11
+ mcm5l1p1_ca_w_0_170_s_0_450 = 1.49e-04  mcm5l1p1_cc_w_0_170_s_0_450 = 3.25e-11  mcm5l1p1_cf_w_0_170_s_0_450 = 2.58e-11
+ mcm5l1p1_ca_w_0_170_s_0_540 = 1.49e-04  mcm5l1p1_cc_w_0_170_s_0_540 = 2.58e-11  mcm5l1p1_cf_w_0_170_s_0_540 = 2.98e-11
+ mcm5l1p1_ca_w_0_170_s_0_720 = 1.49e-04  mcm5l1p1_cc_w_0_170_s_0_720 = 1.76e-11  mcm5l1p1_cf_w_0_170_s_0_720 = 3.55e-11
+ mcm5l1p1_ca_w_0_170_s_1_080 = 1.49e-04  mcm5l1p1_cc_w_0_170_s_1_080 = 9.17e-12  mcm5l1p1_cf_w_0_170_s_1_080 = 4.24e-11
+ mcm5l1p1_ca_w_0_170_s_1_980 = 1.49e-04  mcm5l1p1_cc_w_0_170_s_1_980 = 2.72e-12  mcm5l1p1_cf_w_0_170_s_1_980 = 4.84e-11
+ mcm5l1p1_ca_w_0_170_s_4_500 = 1.49e-04  mcm5l1p1_cc_w_0_170_s_4_500 = 2.88e-13  mcm5l1p1_cf_w_0_170_s_4_500 = 5.08e-11
+ mcm5l1p1_ca_w_1_360_s_0_180 = 1.49e-04  mcm5l1p1_cc_w_1_360_s_0_180 = 9.62e-11  mcm5l1p1_cf_w_1_360_s_0_180 = 1.11e-11
+ mcm5l1p1_ca_w_1_360_s_0_225 = 1.49e-04  mcm5l1p1_cc_w_1_360_s_0_225 = 7.87e-11  mcm5l1p1_cf_w_1_360_s_0_225 = 1.40e-11
+ mcm5l1p1_ca_w_1_360_s_0_270 = 1.49e-04  mcm5l1p1_cc_w_1_360_s_0_270 = 6.69e-11  mcm5l1p1_cf_w_1_360_s_0_270 = 1.67e-11
+ mcm5l1p1_ca_w_1_360_s_0_360 = 1.49e-04  mcm5l1p1_cc_w_1_360_s_0_360 = 5.14e-11  mcm5l1p1_cf_w_1_360_s_0_360 = 2.17e-11
+ mcm5l1p1_ca_w_1_360_s_0_450 = 1.49e-04  mcm5l1p1_cc_w_1_360_s_0_450 = 4.15e-11  mcm5l1p1_cf_w_1_360_s_0_450 = 2.60e-11
+ mcm5l1p1_ca_w_1_360_s_0_540 = 1.49e-04  mcm5l1p1_cc_w_1_360_s_0_540 = 3.45e-11  mcm5l1p1_cf_w_1_360_s_0_540 = 2.98e-11
+ mcm5l1p1_ca_w_1_360_s_0_720 = 1.49e-04  mcm5l1p1_cc_w_1_360_s_0_720 = 2.50e-11  mcm5l1p1_cf_w_1_360_s_0_720 = 3.60e-11
+ mcm5l1p1_ca_w_1_360_s_1_080 = 1.49e-04  mcm5l1p1_cc_w_1_360_s_1_080 = 1.48e-11  mcm5l1p1_cf_w_1_360_s_1_080 = 4.39e-11
+ mcm5l1p1_ca_w_1_360_s_1_980 = 1.49e-04  mcm5l1p1_cc_w_1_360_s_1_980 = 5.31e-12  mcm5l1p1_cf_w_1_360_s_1_980 = 5.24e-11
+ mcm5l1p1_ca_w_1_360_s_4_500 = 1.49e-04  mcm5l1p1_cc_w_1_360_s_4_500 = 6.90e-13  mcm5l1p1_cf_w_1_360_s_4_500 = 5.69e-11
+ mcrdll1f_ca_w_0_170_s_0_180 = 4.87e-05  mcrdll1f_cc_w_0_170_s_0_180 = 9.28e-11  mcrdll1f_cf_w_0_170_s_0_180 = 3.74e-12
+ mcrdll1f_ca_w_0_170_s_0_225 = 4.87e-05  mcrdll1f_cc_w_0_170_s_0_225 = 7.67e-11  mcrdll1f_cf_w_0_170_s_0_225 = 4.79e-12
+ mcrdll1f_ca_w_0_170_s_0_270 = 4.87e-05  mcrdll1f_cc_w_0_170_s_0_270 = 6.65e-11  mcrdll1f_cf_w_0_170_s_0_270 = 5.79e-12
+ mcrdll1f_ca_w_0_170_s_0_360 = 4.87e-05  mcrdll1f_cc_w_0_170_s_0_360 = 5.28e-11  mcrdll1f_cf_w_0_170_s_0_360 = 7.94e-12
+ mcrdll1f_ca_w_0_170_s_0_450 = 4.87e-05  mcrdll1f_cc_w_0_170_s_0_450 = 4.44e-11  mcrdll1f_cf_w_0_170_s_0_450 = 9.66e-12
+ mcrdll1f_ca_w_0_170_s_0_540 = 4.87e-05  mcrdll1f_cc_w_0_170_s_0_540 = 3.81e-11  mcrdll1f_cf_w_0_170_s_0_540 = 1.17e-11
+ mcrdll1f_ca_w_0_170_s_0_720 = 4.87e-05  mcrdll1f_cc_w_0_170_s_0_720 = 2.96e-11  mcrdll1f_cf_w_0_170_s_0_720 = 1.50e-11
+ mcrdll1f_ca_w_0_170_s_1_080 = 4.87e-05  mcrdll1f_cc_w_0_170_s_1_080 = 1.98e-11  mcrdll1f_cf_w_0_170_s_1_080 = 2.05e-11
+ mcrdll1f_ca_w_0_170_s_1_980 = 4.87e-05  mcrdll1f_cc_w_0_170_s_1_980 = 9.18e-12  mcrdll1f_cf_w_0_170_s_1_980 = 2.84e-11
+ mcrdll1f_ca_w_0_170_s_4_500 = 4.87e-05  mcrdll1f_cc_w_0_170_s_4_500 = 1.98e-12  mcrdll1f_cf_w_0_170_s_4_500 = 3.50e-11
+ mcrdll1f_ca_w_1_360_s_0_180 = 4.87e-05  mcrdll1f_cc_w_1_360_s_0_180 = 1.12e-10  mcrdll1f_cf_w_1_360_s_0_180 = 3.74e-12
+ mcrdll1f_ca_w_1_360_s_0_225 = 4.87e-05  mcrdll1f_cc_w_1_360_s_0_225 = 9.43e-11  mcrdll1f_cf_w_1_360_s_0_225 = 4.78e-12
+ mcrdll1f_ca_w_1_360_s_0_270 = 4.87e-05  mcrdll1f_cc_w_1_360_s_0_270 = 8.25e-11  mcrdll1f_cf_w_1_360_s_0_270 = 5.80e-12
+ mcrdll1f_ca_w_1_360_s_0_360 = 4.87e-05  mcrdll1f_cc_w_1_360_s_0_360 = 6.72e-11  mcrdll1f_cf_w_1_360_s_0_360 = 7.81e-12
+ mcrdll1f_ca_w_1_360_s_0_450 = 4.87e-05  mcrdll1f_cc_w_1_360_s_0_450 = 5.72e-11  mcrdll1f_cf_w_1_360_s_0_450 = 9.73e-12
+ mcrdll1f_ca_w_1_360_s_0_540 = 4.87e-05  mcrdll1f_cc_w_1_360_s_0_540 = 5.01e-11  mcrdll1f_cf_w_1_360_s_0_540 = 1.15e-11
+ mcrdll1f_ca_w_1_360_s_0_720 = 4.87e-05  mcrdll1f_cc_w_1_360_s_0_720 = 4.01e-11  mcrdll1f_cf_w_1_360_s_0_720 = 1.49e-11
+ mcrdll1f_ca_w_1_360_s_1_080 = 4.87e-05  mcrdll1f_cc_w_1_360_s_1_080 = 2.84e-11  mcrdll1f_cf_w_1_360_s_1_080 = 2.07e-11
+ mcrdll1f_ca_w_1_360_s_1_980 = 4.87e-05  mcrdll1f_cc_w_1_360_s_1_980 = 1.46e-11  mcrdll1f_cf_w_1_360_s_1_980 = 3.03e-11
+ mcrdll1f_ca_w_1_360_s_4_500 = 4.87e-05  mcrdll1f_cc_w_1_360_s_4_500 = 3.89e-12  mcrdll1f_cf_w_1_360_s_4_500 = 3.98e-11
+ mcrdll1d_ca_w_0_170_s_0_180 = 6.92e-05  mcrdll1d_cc_w_0_170_s_0_180 = 9.06e-11  mcrdll1d_cf_w_0_170_s_0_180 = 5.26e-12
+ mcrdll1d_ca_w_0_170_s_0_225 = 6.92e-05  mcrdll1d_cc_w_0_170_s_0_225 = 7.40e-11  mcrdll1d_cf_w_0_170_s_0_225 = 6.72e-12
+ mcrdll1d_ca_w_0_170_s_0_270 = 6.92e-05  mcrdll1d_cc_w_0_170_s_0_270 = 6.36e-11  mcrdll1d_cf_w_0_170_s_0_270 = 8.10e-12
+ mcrdll1d_ca_w_0_170_s_0_360 = 6.92e-05  mcrdll1d_cc_w_0_170_s_0_360 = 4.97e-11  mcrdll1d_cf_w_0_170_s_0_360 = 1.10e-11
+ mcrdll1d_ca_w_0_170_s_0_450 = 6.92e-05  mcrdll1d_cc_w_0_170_s_0_450 = 4.12e-11  mcrdll1d_cf_w_0_170_s_0_450 = 1.33e-11
+ mcrdll1d_ca_w_0_170_s_0_540 = 6.92e-05  mcrdll1d_cc_w_0_170_s_0_540 = 3.46e-11  mcrdll1d_cf_w_0_170_s_0_540 = 1.59e-11
+ mcrdll1d_ca_w_0_170_s_0_720 = 6.92e-05  mcrdll1d_cc_w_0_170_s_0_720 = 2.61e-11  mcrdll1d_cf_w_0_170_s_0_720 = 2.01e-11
+ mcrdll1d_ca_w_0_170_s_1_080 = 6.92e-05  mcrdll1d_cc_w_0_170_s_1_080 = 1.64e-11  mcrdll1d_cf_w_0_170_s_1_080 = 2.65e-11
+ mcrdll1d_ca_w_0_170_s_1_980 = 6.92e-05  mcrdll1d_cc_w_0_170_s_1_980 = 6.87e-12  mcrdll1d_cf_w_0_170_s_1_980 = 3.44e-11
+ mcrdll1d_ca_w_0_170_s_4_500 = 6.92e-05  mcrdll1d_cc_w_0_170_s_4_500 = 1.35e-12  mcrdll1d_cf_w_0_170_s_4_500 = 3.96e-11
+ mcrdll1d_ca_w_1_360_s_0_180 = 6.92e-05  mcrdll1d_cc_w_1_360_s_0_180 = 1.08e-10  mcrdll1d_cf_w_1_360_s_0_180 = 5.27e-12
+ mcrdll1d_ca_w_1_360_s_0_225 = 6.92e-05  mcrdll1d_cc_w_1_360_s_0_225 = 9.02e-11  mcrdll1d_cf_w_1_360_s_0_225 = 6.71e-12
+ mcrdll1d_ca_w_1_360_s_0_270 = 6.92e-05  mcrdll1d_cc_w_1_360_s_0_270 = 7.84e-11  mcrdll1d_cf_w_1_360_s_0_270 = 8.11e-12
+ mcrdll1d_ca_w_1_360_s_0_360 = 6.92e-05  mcrdll1d_cc_w_1_360_s_0_360 = 6.31e-11  mcrdll1d_cf_w_1_360_s_0_360 = 1.08e-11
+ mcrdll1d_ca_w_1_360_s_0_450 = 6.92e-05  mcrdll1d_cc_w_1_360_s_0_450 = 5.32e-11  mcrdll1d_cf_w_1_360_s_0_450 = 1.34e-11
+ mcrdll1d_ca_w_1_360_s_0_540 = 6.92e-05  mcrdll1d_cc_w_1_360_s_0_540 = 4.60e-11  mcrdll1d_cf_w_1_360_s_0_540 = 1.58e-11
+ mcrdll1d_ca_w_1_360_s_0_720 = 6.92e-05  mcrdll1d_cc_w_1_360_s_0_720 = 3.61e-11  mcrdll1d_cf_w_1_360_s_0_720 = 2.01e-11
+ mcrdll1d_ca_w_1_360_s_1_080 = 6.92e-05  mcrdll1d_cc_w_1_360_s_1_080 = 2.47e-11  mcrdll1d_cf_w_1_360_s_1_080 = 2.69e-11
+ mcrdll1d_ca_w_1_360_s_1_980 = 6.92e-05  mcrdll1d_cc_w_1_360_s_1_980 = 1.19e-11  mcrdll1d_cf_w_1_360_s_1_980 = 3.69e-11
+ mcrdll1d_ca_w_1_360_s_4_500 = 6.92e-05  mcrdll1d_cc_w_1_360_s_4_500 = 2.98e-12  mcrdll1d_cf_w_1_360_s_4_500 = 4.53e-11
+ mcrdll1p1_ca_w_0_170_s_0_180 = 1.44e-04  mcrdll1p1_cc_w_0_170_s_0_180 = 8.38e-11  mcrdll1p1_cf_w_0_170_s_0_180 = 1.06e-11
+ mcrdll1p1_ca_w_0_170_s_0_225 = 1.44e-04  mcrdll1p1_cc_w_0_170_s_0_225 = 6.71e-11  mcrdll1p1_cf_w_0_170_s_0_225 = 1.33e-11
+ mcrdll1p1_ca_w_0_170_s_0_270 = 1.44e-04  mcrdll1p1_cc_w_0_170_s_0_270 = 5.66e-11  mcrdll1p1_cf_w_0_170_s_0_270 = 1.59e-11
+ mcrdll1p1_ca_w_0_170_s_0_360 = 1.44e-04  mcrdll1p1_cc_w_0_170_s_0_360 = 4.22e-11  mcrdll1p1_cf_w_0_170_s_0_360 = 2.10e-11
+ mcrdll1p1_ca_w_0_170_s_0_450 = 1.44e-04  mcrdll1p1_cc_w_0_170_s_0_450 = 3.37e-11  mcrdll1p1_cf_w_0_170_s_0_450 = 2.48e-11
+ mcrdll1p1_ca_w_0_170_s_0_540 = 1.44e-04  mcrdll1p1_cc_w_0_170_s_0_540 = 2.70e-11  mcrdll1p1_cf_w_0_170_s_0_540 = 2.88e-11
+ mcrdll1p1_ca_w_0_170_s_0_720 = 1.44e-04  mcrdll1p1_cc_w_0_170_s_0_720 = 1.89e-11  mcrdll1p1_cf_w_0_170_s_0_720 = 3.44e-11
+ mcrdll1p1_ca_w_0_170_s_1_080 = 1.44e-04  mcrdll1p1_cc_w_0_170_s_1_080 = 1.03e-11  mcrdll1p1_cf_w_0_170_s_1_080 = 4.15e-11
+ mcrdll1p1_ca_w_0_170_s_1_980 = 1.44e-04  mcrdll1p1_cc_w_0_170_s_1_980 = 3.72e-12  mcrdll1p1_cf_w_0_170_s_1_980 = 4.77e-11
+ mcrdll1p1_ca_w_0_170_s_4_500 = 1.44e-04  mcrdll1p1_cc_w_0_170_s_4_500 = 6.76e-13  mcrdll1p1_cf_w_0_170_s_4_500 = 5.06e-11
+ mcrdll1p1_ca_w_1_360_s_0_180 = 1.44e-04  mcrdll1p1_cc_w_1_360_s_0_180 = 9.97e-11  mcrdll1p1_cf_w_1_360_s_0_180 = 1.07e-11
+ mcrdll1p1_ca_w_1_360_s_0_225 = 1.44e-04  mcrdll1p1_cc_w_1_360_s_0_225 = 8.21e-11  mcrdll1p1_cf_w_1_360_s_0_225 = 1.35e-11
+ mcrdll1p1_ca_w_1_360_s_0_270 = 1.44e-04  mcrdll1p1_cc_w_1_360_s_0_270 = 7.04e-11  mcrdll1p1_cf_w_1_360_s_0_270 = 1.61e-11
+ mcrdll1p1_ca_w_1_360_s_0_360 = 1.44e-04  mcrdll1p1_cc_w_1_360_s_0_360 = 5.51e-11  mcrdll1p1_cf_w_1_360_s_0_360 = 2.09e-11
+ mcrdll1p1_ca_w_1_360_s_0_450 = 1.44e-04  mcrdll1p1_cc_w_1_360_s_0_450 = 4.53e-11  mcrdll1p1_cf_w_1_360_s_0_450 = 2.51e-11
+ mcrdll1p1_ca_w_1_360_s_0_540 = 1.44e-04  mcrdll1p1_cc_w_1_360_s_0_540 = 3.83e-11  mcrdll1p1_cf_w_1_360_s_0_540 = 2.88e-11
+ mcrdll1p1_ca_w_1_360_s_0_720 = 1.44e-04  mcrdll1p1_cc_w_1_360_s_0_720 = 2.89e-11  mcrdll1p1_cf_w_1_360_s_0_720 = 3.48e-11
+ mcrdll1p1_ca_w_1_360_s_1_080 = 1.44e-04  mcrdll1p1_cc_w_1_360_s_1_080 = 1.85e-11  mcrdll1p1_cf_w_1_360_s_1_080 = 4.29e-11
+ mcrdll1p1_ca_w_1_360_s_1_980 = 1.44e-04  mcrdll1p1_cc_w_1_360_s_1_980 = 8.24e-12  mcrdll1p1_cf_w_1_360_s_1_980 = 5.21e-11
+ mcrdll1p1_ca_w_1_360_s_4_500 = 1.44e-04  mcrdll1p1_cc_w_1_360_s_4_500 = 1.98e-12  mcrdll1p1_cf_w_1_360_s_4_500 = 5.81e-11
+ mcm2m1f_ca_w_0_140_s_0_140 = 2.50e-04  mcm2m1f_cc_w_0_140_s_0_140 = 1.03e-10  mcm2m1f_cf_w_0_140_s_0_140 = 1.29e-11
+ mcm2m1f_ca_w_0_140_s_0_175 = 2.50e-04  mcm2m1f_cc_w_0_140_s_0_175 = 9.85e-11  mcm2m1f_cf_w_0_140_s_0_175 = 1.63e-11
+ mcm2m1f_ca_w_0_140_s_0_210 = 2.50e-04  mcm2m1f_cc_w_0_140_s_0_210 = 9.18e-11  mcm2m1f_cf_w_0_140_s_0_210 = 1.94e-11
+ mcm2m1f_ca_w_0_140_s_0_280 = 2.50e-04  mcm2m1f_cc_w_0_140_s_0_280 = 7.51e-11  mcm2m1f_cf_w_0_140_s_0_280 = 2.52e-11
+ mcm2m1f_ca_w_0_140_s_0_350 = 2.50e-04  mcm2m1f_cc_w_0_140_s_0_350 = 6.07e-11  mcm2m1f_cf_w_0_140_s_0_350 = 3.05e-11
+ mcm2m1f_ca_w_0_140_s_0_420 = 2.50e-04  mcm2m1f_cc_w_0_140_s_0_420 = 4.92e-11  mcm2m1f_cf_w_0_140_s_0_420 = 3.54e-11
+ mcm2m1f_ca_w_0_140_s_0_560 = 2.50e-04  mcm2m1f_cc_w_0_140_s_0_560 = 3.35e-11  mcm2m1f_cf_w_0_140_s_0_560 = 4.30e-11
+ mcm2m1f_ca_w_0_140_s_0_840 = 2.50e-04  mcm2m1f_cc_w_0_140_s_0_840 = 1.75e-11  mcm2m1f_cf_w_0_140_s_0_840 = 5.39e-11
+ mcm2m1f_ca_w_0_140_s_1_540 = 2.50e-04  mcm2m1f_cc_w_0_140_s_1_540 = 4.32e-12  mcm2m1f_cf_w_0_140_s_1_540 = 6.54e-11
+ mcm2m1f_ca_w_0_140_s_3_500 = 2.50e-04  mcm2m1f_cc_w_0_140_s_3_500 = 1.95e-13  mcm2m1f_cf_w_0_140_s_3_500 = 7.00e-11
+ mcm2m1f_ca_w_1_120_s_0_140 = 2.50e-04  mcm2m1f_cc_w_1_120_s_0_140 = 1.11e-10  mcm2m1f_cf_w_1_120_s_0_140 = 1.29e-11
+ mcm2m1f_ca_w_1_120_s_0_175 = 2.50e-04  mcm2m1f_cc_w_1_120_s_0_175 = 1.06e-10  mcm2m1f_cf_w_1_120_s_0_175 = 1.63e-11
+ mcm2m1f_ca_w_1_120_s_0_210 = 2.50e-04  mcm2m1f_cc_w_1_120_s_0_210 = 9.83e-11  mcm2m1f_cf_w_1_120_s_0_210 = 1.94e-11
+ mcm2m1f_ca_w_1_120_s_0_280 = 2.50e-04  mcm2m1f_cc_w_1_120_s_0_280 = 8.04e-11  mcm2m1f_cf_w_1_120_s_0_280 = 2.52e-11
+ mcm2m1f_ca_w_1_120_s_0_350 = 2.50e-04  mcm2m1f_cc_w_1_120_s_0_350 = 6.55e-11  mcm2m1f_cf_w_1_120_s_0_350 = 3.05e-11
+ mcm2m1f_ca_w_1_120_s_0_420 = 2.50e-04  mcm2m1f_cc_w_1_120_s_0_420 = 5.31e-11  mcm2m1f_cf_w_1_120_s_0_420 = 3.53e-11
+ mcm2m1f_ca_w_1_120_s_0_560 = 2.50e-04  mcm2m1f_cc_w_1_120_s_0_560 = 3.63e-11  mcm2m1f_cf_w_1_120_s_0_560 = 4.31e-11
+ mcm2m1f_ca_w_1_120_s_0_840 = 2.50e-04  mcm2m1f_cc_w_1_120_s_0_840 = 1.92e-11  mcm2m1f_cf_w_1_120_s_0_840 = 5.42e-11
+ mcm2m1f_ca_w_1_120_s_1_540 = 2.50e-04  mcm2m1f_cc_w_1_120_s_1_540 = 4.95e-12  mcm2m1f_cf_w_1_120_s_1_540 = 6.65e-11
+ mcm2m1f_ca_w_1_120_s_3_500 = 2.50e-04  mcm2m1f_cc_w_1_120_s_3_500 = 2.05e-13  mcm2m1f_cf_w_1_120_s_3_500 = 7.13e-11
+ mcm2m1d_ca_w_0_140_s_0_140 = 2.59e-04  mcm2m1d_cc_w_0_140_s_0_140 = 1.03e-10  mcm2m1d_cf_w_0_140_s_0_140 = 1.34e-11
+ mcm2m1d_ca_w_0_140_s_0_175 = 2.59e-04  mcm2m1d_cc_w_0_140_s_0_175 = 9.73e-11  mcm2m1d_cf_w_0_140_s_0_175 = 1.70e-11
+ mcm2m1d_ca_w_0_140_s_0_210 = 2.59e-04  mcm2m1d_cc_w_0_140_s_0_210 = 9.04e-11  mcm2m1d_cf_w_0_140_s_0_210 = 2.02e-11
+ mcm2m1d_ca_w_0_140_s_0_280 = 2.59e-04  mcm2m1d_cc_w_0_140_s_0_280 = 7.36e-11  mcm2m1d_cf_w_0_140_s_0_280 = 2.63e-11
+ mcm2m1d_ca_w_0_140_s_0_350 = 2.59e-04  mcm2m1d_cc_w_0_140_s_0_350 = 5.97e-11  mcm2m1d_cf_w_0_140_s_0_350 = 3.18e-11
+ mcm2m1d_ca_w_0_140_s_0_420 = 2.59e-04  mcm2m1d_cc_w_0_140_s_0_420 = 4.75e-11  mcm2m1d_cf_w_0_140_s_0_420 = 3.70e-11
+ mcm2m1d_ca_w_0_140_s_0_560 = 2.59e-04  mcm2m1d_cc_w_0_140_s_0_560 = 3.17e-11  mcm2m1d_cf_w_0_140_s_0_560 = 4.51e-11
+ mcm2m1d_ca_w_0_140_s_0_840 = 2.59e-04  mcm2m1d_cc_w_0_140_s_0_840 = 1.56e-11  mcm2m1d_cf_w_0_140_s_0_840 = 5.63e-11
+ mcm2m1d_ca_w_0_140_s_1_540 = 2.59e-04  mcm2m1d_cc_w_0_140_s_1_540 = 3.32e-12  mcm2m1d_cf_w_0_140_s_1_540 = 6.74e-11
+ mcm2m1d_ca_w_0_140_s_3_500 = 2.59e-04  mcm2m1d_cc_w_0_140_s_3_500 = 1.05e-13  mcm2m1d_cf_w_0_140_s_3_500 = 7.10e-11
+ mcm2m1d_ca_w_1_120_s_0_140 = 2.59e-04  mcm2m1d_cc_w_1_120_s_0_140 = 1.08e-10  mcm2m1d_cf_w_1_120_s_0_140 = 1.35e-11
+ mcm2m1d_ca_w_1_120_s_0_175 = 2.59e-04  mcm2m1d_cc_w_1_120_s_0_175 = 1.03e-10  mcm2m1d_cf_w_1_120_s_0_175 = 1.70e-11
+ mcm2m1d_ca_w_1_120_s_0_210 = 2.59e-04  mcm2m1d_cc_w_1_120_s_0_210 = 9.55e-11  mcm2m1d_cf_w_1_120_s_0_210 = 2.03e-11
+ mcm2m1d_ca_w_1_120_s_0_280 = 2.59e-04  mcm2m1d_cc_w_1_120_s_0_280 = 7.79e-11  mcm2m1d_cf_w_1_120_s_0_280 = 2.64e-11
+ mcm2m1d_ca_w_1_120_s_0_350 = 2.59e-04  mcm2m1d_cc_w_1_120_s_0_350 = 6.30e-11  mcm2m1d_cf_w_1_120_s_0_350 = 3.19e-11
+ mcm2m1d_ca_w_1_120_s_0_420 = 2.59e-04  mcm2m1d_cc_w_1_120_s_0_420 = 5.04e-11  mcm2m1d_cf_w_1_120_s_0_420 = 3.70e-11
+ mcm2m1d_ca_w_1_120_s_0_560 = 2.59e-04  mcm2m1d_cc_w_1_120_s_0_560 = 3.37e-11  mcm2m1d_cf_w_1_120_s_0_560 = 4.53e-11
+ mcm2m1d_ca_w_1_120_s_0_840 = 2.59e-04  mcm2m1d_cc_w_1_120_s_0_840 = 1.68e-11  mcm2m1d_cf_w_1_120_s_0_840 = 5.66e-11
+ mcm2m1d_ca_w_1_120_s_1_540 = 2.59e-04  mcm2m1d_cc_w_1_120_s_1_540 = 3.59e-12  mcm2m1d_cf_w_1_120_s_1_540 = 6.82e-11
+ mcm2m1d_ca_w_1_120_s_3_500 = 2.59e-04  mcm2m1d_cc_w_1_120_s_3_500 = 1.30e-13  mcm2m1d_cf_w_1_120_s_3_500 = 7.21e-11
+ mcm2m1p1_ca_w_0_140_s_0_140 = 2.79e-04  mcm2m1p1_cc_w_0_140_s_0_140 = 1.01e-10  mcm2m1p1_cf_w_0_140_s_0_140 = 1.46e-11
+ mcm2m1p1_ca_w_0_140_s_0_175 = 2.79e-04  mcm2m1p1_cc_w_0_140_s_0_175 = 9.46e-11  mcm2m1p1_cf_w_0_140_s_0_175 = 1.84e-11
+ mcm2m1p1_ca_w_0_140_s_0_210 = 2.79e-04  mcm2m1p1_cc_w_0_140_s_0_210 = 8.80e-11  mcm2m1p1_cf_w_0_140_s_0_210 = 2.21e-11
+ mcm2m1p1_ca_w_0_140_s_0_280 = 2.79e-04  mcm2m1p1_cc_w_0_140_s_0_280 = 7.06e-11  mcm2m1p1_cf_w_0_140_s_0_280 = 2.88e-11
+ mcm2m1p1_ca_w_0_140_s_0_350 = 2.79e-04  mcm2m1p1_cc_w_0_140_s_0_350 = 5.64e-11  mcm2m1p1_cf_w_0_140_s_0_350 = 3.49e-11
+ mcm2m1p1_ca_w_0_140_s_0_420 = 2.79e-04  mcm2m1p1_cc_w_0_140_s_0_420 = 4.40e-11  mcm2m1p1_cf_w_0_140_s_0_420 = 4.05e-11
+ mcm2m1p1_ca_w_0_140_s_0_560 = 2.79e-04  mcm2m1p1_cc_w_0_140_s_0_560 = 2.81e-11  mcm2m1p1_cf_w_0_140_s_0_560 = 4.95e-11
+ mcm2m1p1_ca_w_0_140_s_0_840 = 2.79e-04  mcm2m1p1_cc_w_0_140_s_0_840 = 1.24e-11  mcm2m1p1_cf_w_0_140_s_0_840 = 6.12e-11
+ mcm2m1p1_ca_w_0_140_s_1_540 = 2.79e-04  mcm2m1p1_cc_w_0_140_s_1_540 = 1.86e-12  mcm2m1p1_cf_w_0_140_s_1_540 = 7.14e-11
+ mcm2m1p1_ca_w_0_140_s_3_500 = 2.79e-04  mcm2m1p1_cc_w_0_140_s_3_500 = 3.00e-14  mcm2m1p1_cf_w_0_140_s_3_500 = 7.38e-11
+ mcm2m1p1_ca_w_1_120_s_0_140 = 2.79e-04  mcm2m1p1_cc_w_1_120_s_0_140 = 1.03e-10  mcm2m1p1_cf_w_1_120_s_0_140 = 1.47e-11
+ mcm2m1p1_ca_w_1_120_s_0_175 = 2.79e-04  mcm2m1p1_cc_w_1_120_s_0_175 = 9.80e-11  mcm2m1p1_cf_w_1_120_s_0_175 = 1.86e-11
+ mcm2m1p1_ca_w_1_120_s_0_210 = 2.79e-04  mcm2m1p1_cc_w_1_120_s_0_210 = 9.06e-11  mcm2m1p1_cf_w_1_120_s_0_210 = 2.22e-11
+ mcm2m1p1_ca_w_1_120_s_0_280 = 2.79e-04  mcm2m1p1_cc_w_1_120_s_0_280 = 7.31e-11  mcm2m1p1_cf_w_1_120_s_0_280 = 2.89e-11
+ mcm2m1p1_ca_w_1_120_s_0_350 = 2.79e-04  mcm2m1p1_cc_w_1_120_s_0_350 = 5.79e-11  mcm2m1p1_cf_w_1_120_s_0_350 = 3.50e-11
+ mcm2m1p1_ca_w_1_120_s_0_420 = 2.79e-04  mcm2m1p1_cc_w_1_120_s_0_420 = 4.56e-11  mcm2m1p1_cf_w_1_120_s_0_420 = 4.06e-11
+ mcm2m1p1_ca_w_1_120_s_0_560 = 2.79e-04  mcm2m1p1_cc_w_1_120_s_0_560 = 2.90e-11  mcm2m1p1_cf_w_1_120_s_0_560 = 4.96e-11
+ mcm2m1p1_ca_w_1_120_s_0_840 = 2.79e-04  mcm2m1p1_cc_w_1_120_s_0_840 = 1.29e-11  mcm2m1p1_cf_w_1_120_s_0_840 = 6.16e-11
+ mcm2m1p1_ca_w_1_120_s_1_540 = 2.79e-04  mcm2m1p1_cc_w_1_120_s_1_540 = 1.95e-12  mcm2m1p1_cf_w_1_120_s_1_540 = 7.19e-11
+ mcm2m1p1_ca_w_1_120_s_3_500 = 2.79e-04  mcm2m1p1_cc_w_1_120_s_3_500 = 1.00e-13  mcm2m1p1_cf_w_1_120_s_3_500 = 7.43e-11
+ mcm2m1l1_ca_w_0_140_s_0_140 = 3.81e-04  mcm2m1l1_cc_w_0_140_s_0_140 = 9.17e-11  mcm2m1l1_cf_w_0_140_s_0_140 = 1.99e-11
+ mcm2m1l1_ca_w_0_140_s_0_175 = 3.81e-04  mcm2m1l1_cc_w_0_140_s_0_175 = 8.63e-11  mcm2m1l1_cf_w_0_140_s_0_175 = 2.55e-11
+ mcm2m1l1_ca_w_0_140_s_0_210 = 3.81e-04  mcm2m1l1_cc_w_0_140_s_0_210 = 7.83e-11  mcm2m1l1_cf_w_0_140_s_0_210 = 3.08e-11
+ mcm2m1l1_ca_w_0_140_s_0_280 = 3.81e-04  mcm2m1l1_cc_w_0_140_s_0_280 = 6.15e-11  mcm2m1l1_cf_w_0_140_s_0_280 = 4.04e-11
+ mcm2m1l1_ca_w_0_140_s_0_350 = 3.81e-04  mcm2m1l1_cc_w_0_140_s_0_350 = 4.63e-11  mcm2m1l1_cf_w_0_140_s_0_350 = 4.90e-11
+ mcm2m1l1_ca_w_0_140_s_0_420 = 3.81e-04  mcm2m1l1_cc_w_0_140_s_0_420 = 3.43e-11  mcm2m1l1_cf_w_0_140_s_0_420 = 5.65e-11
+ mcm2m1l1_ca_w_0_140_s_0_560 = 3.81e-04  mcm2m1l1_cc_w_0_140_s_0_560 = 1.90e-11  mcm2m1l1_cf_w_0_140_s_0_560 = 6.79e-11
+ mcm2m1l1_ca_w_0_140_s_0_840 = 3.81e-04  mcm2m1l1_cc_w_0_140_s_0_840 = 6.10e-12  mcm2m1l1_cf_w_0_140_s_0_840 = 8.01e-11
+ mcm2m1l1_ca_w_0_140_s_1_540 = 3.81e-04  mcm2m1l1_cc_w_0_140_s_1_540 = 5.00e-13  mcm2m1l1_cf_w_0_140_s_1_540 = 8.69e-11
+ mcm2m1l1_ca_w_0_140_s_3_500 = 3.81e-04  mcm2m1l1_cc_w_0_140_s_3_500 = 5.00e-14  mcm2m1l1_cf_w_0_140_s_3_500 = 8.81e-11
+ mcm2m1l1_ca_w_1_120_s_0_140 = 3.81e-04  mcm2m1l1_cc_w_1_120_s_0_140 = 9.31e-11  mcm2m1l1_cf_w_1_120_s_0_140 = 2.00e-11
+ mcm2m1l1_ca_w_1_120_s_0_175 = 3.81e-04  mcm2m1l1_cc_w_1_120_s_0_175 = 8.66e-11  mcm2m1l1_cf_w_1_120_s_0_175 = 2.56e-11
+ mcm2m1l1_ca_w_1_120_s_0_210 = 3.81e-04  mcm2m1l1_cc_w_1_120_s_0_210 = 7.91e-11  mcm2m1l1_cf_w_1_120_s_0_210 = 3.09e-11
+ mcm2m1l1_ca_w_1_120_s_0_280 = 3.81e-04  mcm2m1l1_cc_w_1_120_s_0_280 = 6.16e-11  mcm2m1l1_cf_w_1_120_s_0_280 = 4.05e-11
+ mcm2m1l1_ca_w_1_120_s_0_350 = 3.81e-04  mcm2m1l1_cc_w_1_120_s_0_350 = 4.66e-11  mcm2m1l1_cf_w_1_120_s_0_350 = 4.91e-11
+ mcm2m1l1_ca_w_1_120_s_0_420 = 3.81e-04  mcm2m1l1_cc_w_1_120_s_0_420 = 3.45e-11  mcm2m1l1_cf_w_1_120_s_0_420 = 5.67e-11
+ mcm2m1l1_ca_w_1_120_s_0_560 = 3.81e-04  mcm2m1l1_cc_w_1_120_s_0_560 = 1.91e-11  mcm2m1l1_cf_w_1_120_s_0_560 = 6.81e-11
+ mcm2m1l1_ca_w_1_120_s_0_840 = 3.81e-04  mcm2m1l1_cc_w_1_120_s_0_840 = 6.15e-12  mcm2m1l1_cf_w_1_120_s_0_840 = 8.01e-11
+ mcm2m1l1_ca_w_1_120_s_1_540 = 3.81e-04  mcm2m1l1_cc_w_1_120_s_1_540 = 4.50e-13  mcm2m1l1_cf_w_1_120_s_1_540 = 8.70e-11
+ mcm2m1l1_ca_w_1_120_s_3_500 = 3.81e-04  mcm2m1l1_cc_w_1_120_s_3_500 = 5.00e-14  mcm2m1l1_cf_w_1_120_s_3_500 = 8.83e-11
+ mcm3m1f_ca_w_0_140_s_0_140 = 7.26e-05  mcm3m1f_cc_w_0_140_s_0_140 = 1.17e-10  mcm3m1f_cf_w_0_140_s_0_140 = 4.22e-12
+ mcm3m1f_ca_w_0_140_s_0_175 = 7.26e-05  mcm3m1f_cc_w_0_140_s_0_175 = 1.12e-10  mcm3m1f_cf_w_0_140_s_0_175 = 5.44e-12
+ mcm3m1f_ca_w_0_140_s_0_210 = 7.26e-05  mcm3m1f_cc_w_0_140_s_0_210 = 1.06e-10  mcm3m1f_cf_w_0_140_s_0_210 = 6.66e-12
+ mcm3m1f_ca_w_0_140_s_0_280 = 7.26e-05  mcm3m1f_cc_w_0_140_s_0_280 = 9.00e-11  mcm3m1f_cf_w_0_140_s_0_280 = 9.04e-12
+ mcm3m1f_ca_w_0_140_s_0_350 = 7.26e-05  mcm3m1f_cc_w_0_140_s_0_350 = 7.53e-11  mcm3m1f_cf_w_0_140_s_0_350 = 1.14e-11
+ mcm3m1f_ca_w_0_140_s_0_420 = 7.26e-05  mcm3m1f_cc_w_0_140_s_0_420 = 6.32e-11  mcm3m1f_cf_w_0_140_s_0_420 = 1.37e-11
+ mcm3m1f_ca_w_0_140_s_0_560 = 7.26e-05  mcm3m1f_cc_w_0_140_s_0_560 = 4.71e-11  mcm3m1f_cf_w_0_140_s_0_560 = 1.79e-11
+ mcm3m1f_ca_w_0_140_s_0_840 = 7.26e-05  mcm3m1f_cc_w_0_140_s_0_840 = 2.93e-11  mcm3m1f_cf_w_0_140_s_0_840 = 2.53e-11
+ mcm3m1f_ca_w_0_140_s_1_540 = 7.26e-05  mcm3m1f_cc_w_0_140_s_1_540 = 1.07e-11  mcm3m1f_cf_w_0_140_s_1_540 = 3.75e-11
+ mcm3m1f_ca_w_0_140_s_3_500 = 7.26e-05  mcm3m1f_cc_w_0_140_s_3_500 = 8.70e-13  mcm3m1f_cf_w_0_140_s_3_500 = 4.64e-11
+ mcm3m1f_ca_w_1_120_s_0_140 = 7.26e-05  mcm3m1f_cc_w_1_120_s_0_140 = 1.30e-10  mcm3m1f_cf_w_1_120_s_0_140 = 4.26e-12
+ mcm3m1f_ca_w_1_120_s_0_175 = 7.26e-05  mcm3m1f_cc_w_1_120_s_0_175 = 1.24e-10  mcm3m1f_cf_w_1_120_s_0_175 = 5.49e-12
+ mcm3m1f_ca_w_1_120_s_0_210 = 7.26e-05  mcm3m1f_cc_w_1_120_s_0_210 = 1.16e-10  mcm3m1f_cf_w_1_120_s_0_210 = 6.71e-12
+ mcm3m1f_ca_w_1_120_s_0_280 = 7.26e-05  mcm3m1f_cc_w_1_120_s_0_280 = 9.77e-11  mcm3m1f_cf_w_1_120_s_0_280 = 9.11e-12
+ mcm3m1f_ca_w_1_120_s_0_350 = 7.26e-05  mcm3m1f_cc_w_1_120_s_0_350 = 8.21e-11  mcm3m1f_cf_w_1_120_s_0_350 = 1.14e-11
+ mcm3m1f_ca_w_1_120_s_0_420 = 7.26e-05  mcm3m1f_cc_w_1_120_s_0_420 = 6.97e-11  mcm3m1f_cf_w_1_120_s_0_420 = 1.37e-11
+ mcm3m1f_ca_w_1_120_s_0_560 = 7.26e-05  mcm3m1f_cc_w_1_120_s_0_560 = 5.16e-11  mcm3m1f_cf_w_1_120_s_0_560 = 1.80e-11
+ mcm3m1f_ca_w_1_120_s_0_840 = 7.26e-05  mcm3m1f_cc_w_1_120_s_0_840 = 3.21e-11  mcm3m1f_cf_w_1_120_s_0_840 = 2.56e-11
+ mcm3m1f_ca_w_1_120_s_1_540 = 7.26e-05  mcm3m1f_cc_w_1_120_s_1_540 = 1.19e-11  mcm3m1f_cf_w_1_120_s_1_540 = 3.84e-11
+ mcm3m1f_ca_w_1_120_s_3_500 = 7.26e-05  mcm3m1f_cc_w_1_120_s_3_500 = 9.25e-13  mcm3m1f_cf_w_1_120_s_3_500 = 4.82e-11
+ mcm3m1d_ca_w_0_140_s_0_140 = 8.16e-05  mcm3m1d_cc_w_0_140_s_0_140 = 1.15e-10  mcm3m1d_cf_w_0_140_s_0_140 = 4.74e-12
+ mcm3m1d_ca_w_0_140_s_0_175 = 8.16e-05  mcm3m1d_cc_w_0_140_s_0_175 = 1.11e-10  mcm3m1d_cf_w_0_140_s_0_175 = 6.11e-12
+ mcm3m1d_ca_w_0_140_s_0_210 = 8.16e-05  mcm3m1d_cc_w_0_140_s_0_210 = 1.04e-10  mcm3m1d_cf_w_0_140_s_0_210 = 7.49e-12
+ mcm3m1d_ca_w_0_140_s_0_280 = 8.16e-05  mcm3m1d_cc_w_0_140_s_0_280 = 8.85e-11  mcm3m1d_cf_w_0_140_s_0_280 = 1.02e-11
+ mcm3m1d_ca_w_0_140_s_0_350 = 8.16e-05  mcm3m1d_cc_w_0_140_s_0_350 = 7.37e-11  mcm3m1d_cf_w_0_140_s_0_350 = 1.28e-11
+ mcm3m1d_ca_w_0_140_s_0_420 = 8.16e-05  mcm3m1d_cc_w_0_140_s_0_420 = 6.20e-11  mcm3m1d_cf_w_0_140_s_0_420 = 1.53e-11
+ mcm3m1d_ca_w_0_140_s_0_560 = 8.16e-05  mcm3m1d_cc_w_0_140_s_0_560 = 4.52e-11  mcm3m1d_cf_w_0_140_s_0_560 = 2.00e-11
+ mcm3m1d_ca_w_0_140_s_0_840 = 8.16e-05  mcm3m1d_cc_w_0_140_s_0_840 = 2.72e-11  mcm3m1d_cf_w_0_140_s_0_840 = 2.81e-11
+ mcm3m1d_ca_w_0_140_s_1_540 = 8.16e-05  mcm3m1d_cc_w_0_140_s_1_540 = 9.11e-12  mcm3m1d_cf_w_0_140_s_1_540 = 4.06e-11
+ mcm3m1d_ca_w_0_140_s_3_500 = 8.16e-05  mcm3m1d_cc_w_0_140_s_3_500 = 5.80e-13  mcm3m1d_cf_w_0_140_s_3_500 = 4.87e-11
+ mcm3m1d_ca_w_1_120_s_0_140 = 8.16e-05  mcm3m1d_cc_w_1_120_s_0_140 = 1.27e-10  mcm3m1d_cf_w_1_120_s_0_140 = 4.79e-12
+ mcm3m1d_ca_w_1_120_s_0_175 = 8.16e-05  mcm3m1d_cc_w_1_120_s_0_175 = 1.21e-10  mcm3m1d_cf_w_1_120_s_0_175 = 6.18e-12
+ mcm3m1d_ca_w_1_120_s_0_210 = 8.16e-05  mcm3m1d_cc_w_1_120_s_0_210 = 1.13e-10  mcm3m1d_cf_w_1_120_s_0_210 = 7.55e-12
+ mcm3m1d_ca_w_1_120_s_0_280 = 8.16e-05  mcm3m1d_cc_w_1_120_s_0_280 = 9.49e-11  mcm3m1d_cf_w_1_120_s_0_280 = 1.02e-11
+ mcm3m1d_ca_w_1_120_s_0_350 = 8.16e-05  mcm3m1d_cc_w_1_120_s_0_350 = 7.92e-11  mcm3m1d_cf_w_1_120_s_0_350 = 1.29e-11
+ mcm3m1d_ca_w_1_120_s_0_420 = 8.16e-05  mcm3m1d_cc_w_1_120_s_0_420 = 6.66e-11  mcm3m1d_cf_w_1_120_s_0_420 = 1.54e-11
+ mcm3m1d_ca_w_1_120_s_0_560 = 8.16e-05  mcm3m1d_cc_w_1_120_s_0_560 = 4.88e-11  mcm3m1d_cf_w_1_120_s_0_560 = 2.02e-11
+ mcm3m1d_ca_w_1_120_s_0_840 = 8.16e-05  mcm3m1d_cc_w_1_120_s_0_840 = 2.94e-11  mcm3m1d_cf_w_1_120_s_0_840 = 2.84e-11
+ mcm3m1d_ca_w_1_120_s_1_540 = 8.16e-05  mcm3m1d_cc_w_1_120_s_1_540 = 9.94e-12  mcm3m1d_cf_w_1_120_s_1_540 = 4.17e-11
+ mcm3m1d_ca_w_1_120_s_3_500 = 8.16e-05  mcm3m1d_cc_w_1_120_s_3_500 = 5.95e-13  mcm3m1d_cf_w_1_120_s_3_500 = 5.02e-11
+ mcm3m1p1_ca_w_0_140_s_0_140 = 1.02e-04  mcm3m1p1_cc_w_0_140_s_0_140 = 1.12e-10  mcm3m1p1_cf_w_0_140_s_0_140 = 5.90e-12
+ mcm3m1p1_ca_w_0_140_s_0_175 = 1.02e-04  mcm3m1p1_cc_w_0_140_s_0_175 = 1.08e-10  mcm3m1p1_cf_w_0_140_s_0_175 = 7.62e-12
+ mcm3m1p1_ca_w_0_140_s_0_210 = 1.02e-04  mcm3m1p1_cc_w_0_140_s_0_210 = 1.02e-10  mcm3m1p1_cf_w_0_140_s_0_210 = 9.33e-12
+ mcm3m1p1_ca_w_0_140_s_0_280 = 1.02e-04  mcm3m1p1_cc_w_0_140_s_0_280 = 8.56e-11  mcm3m1p1_cf_w_0_140_s_0_280 = 1.27e-11
+ mcm3m1p1_ca_w_0_140_s_0_350 = 1.02e-04  mcm3m1p1_cc_w_0_140_s_0_350 = 7.05e-11  mcm3m1p1_cf_w_0_140_s_0_350 = 1.59e-11
+ mcm3m1p1_ca_w_0_140_s_0_420 = 1.02e-04  mcm3m1p1_cc_w_0_140_s_0_420 = 5.85e-11  mcm3m1p1_cf_w_0_140_s_0_420 = 1.90e-11
+ mcm3m1p1_ca_w_0_140_s_0_560 = 1.02e-04  mcm3m1p1_cc_w_0_140_s_0_560 = 4.15e-11  mcm3m1p1_cf_w_0_140_s_0_560 = 2.46e-11
+ mcm3m1p1_ca_w_0_140_s_0_840 = 1.02e-04  mcm3m1p1_cc_w_0_140_s_0_840 = 2.35e-11  mcm3m1p1_cf_w_0_140_s_0_840 = 3.39e-11
+ mcm3m1p1_ca_w_0_140_s_1_540 = 1.02e-04  mcm3m1p1_cc_w_0_140_s_1_540 = 6.72e-12  mcm3m1p1_cf_w_0_140_s_1_540 = 4.68e-11
+ mcm3m1p1_ca_w_0_140_s_3_500 = 1.02e-04  mcm3m1p1_cc_w_0_140_s_3_500 = 3.05e-13  mcm3m1p1_cf_w_0_140_s_3_500 = 5.31e-11
+ mcm3m1p1_ca_w_1_120_s_0_140 = 1.02e-04  mcm3m1p1_cc_w_1_120_s_0_140 = 1.23e-10  mcm3m1p1_cf_w_1_120_s_0_140 = 6.06e-12
+ mcm3m1p1_ca_w_1_120_s_0_175 = 1.02e-04  mcm3m1p1_cc_w_1_120_s_0_175 = 1.16e-10  mcm3m1p1_cf_w_1_120_s_0_175 = 7.79e-12
+ mcm3m1p1_ca_w_1_120_s_0_210 = 1.02e-04  mcm3m1p1_cc_w_1_120_s_0_210 = 1.08e-10  mcm3m1p1_cf_w_1_120_s_0_210 = 9.49e-12
+ mcm3m1p1_ca_w_1_120_s_0_280 = 1.02e-04  mcm3m1p1_cc_w_1_120_s_0_280 = 9.00e-11  mcm3m1p1_cf_w_1_120_s_0_280 = 1.28e-11
+ mcm3m1p1_ca_w_1_120_s_0_350 = 1.02e-04  mcm3m1p1_cc_w_1_120_s_0_350 = 7.45e-11  mcm3m1p1_cf_w_1_120_s_0_350 = 1.60e-11
+ mcm3m1p1_ca_w_1_120_s_0_420 = 1.02e-04  mcm3m1p1_cc_w_1_120_s_0_420 = 6.21e-11  mcm3m1p1_cf_w_1_120_s_0_420 = 1.91e-11
+ mcm3m1p1_ca_w_1_120_s_0_560 = 1.02e-04  mcm3m1p1_cc_w_1_120_s_0_560 = 4.43e-11  mcm3m1p1_cf_w_1_120_s_0_560 = 2.48e-11
+ mcm3m1p1_ca_w_1_120_s_0_840 = 1.02e-04  mcm3m1p1_cc_w_1_120_s_0_840 = 2.50e-11  mcm3m1p1_cf_w_1_120_s_0_840 = 3.43e-11
+ mcm3m1p1_ca_w_1_120_s_1_540 = 1.02e-04  mcm3m1p1_cc_w_1_120_s_1_540 = 7.17e-12  mcm3m1p1_cf_w_1_120_s_1_540 = 4.77e-11
+ mcm3m1p1_ca_w_1_120_s_3_500 = 1.02e-04  mcm3m1p1_cc_w_1_120_s_3_500 = 3.25e-13  mcm3m1p1_cf_w_1_120_s_3_500 = 5.46e-11
+ mcm3m1l1_ca_w_0_140_s_0_140 = 2.04e-04  mcm3m1l1_cc_w_0_140_s_0_140 = 1.06e-10  mcm3m1l1_cf_w_0_140_s_0_140 = 1.12e-11
+ mcm3m1l1_ca_w_0_140_s_0_175 = 2.04e-04  mcm3m1l1_cc_w_0_140_s_0_175 = 9.96e-11  mcm3m1l1_cf_w_0_140_s_0_175 = 1.47e-11
+ mcm3m1l1_ca_w_0_140_s_0_210 = 2.04e-04  mcm3m1l1_cc_w_0_140_s_0_210 = 9.16e-11  mcm3m1l1_cf_w_0_140_s_0_210 = 1.80e-11
+ mcm3m1l1_ca_w_0_140_s_0_280 = 2.04e-04  mcm3m1l1_cc_w_0_140_s_0_280 = 7.55e-11  mcm3m1l1_cf_w_0_140_s_0_280 = 2.43e-11
+ mcm3m1l1_ca_w_0_140_s_0_350 = 2.04e-04  mcm3m1l1_cc_w_0_140_s_0_350 = 6.06e-11  mcm3m1l1_cf_w_0_140_s_0_350 = 2.99e-11
+ mcm3m1l1_ca_w_0_140_s_0_420 = 2.04e-04  mcm3m1l1_cc_w_0_140_s_0_420 = 4.84e-11  mcm3m1l1_cf_w_0_140_s_0_420 = 3.52e-11
+ mcm3m1l1_ca_w_0_140_s_0_560 = 2.04e-04  mcm3m1l1_cc_w_0_140_s_0_560 = 3.22e-11  mcm3m1l1_cf_w_0_140_s_0_560 = 4.39e-11
+ mcm3m1l1_ca_w_0_140_s_0_840 = 2.04e-04  mcm3m1l1_cc_w_0_140_s_0_840 = 1.56e-11  mcm3m1l1_cf_w_0_140_s_0_840 = 5.57e-11
+ mcm3m1l1_ca_w_0_140_s_1_540 = 2.04e-04  mcm3m1l1_cc_w_0_140_s_1_540 = 3.10e-12  mcm3m1l1_cf_w_0_140_s_1_540 = 6.74e-11
+ mcm3m1l1_ca_w_0_140_s_3_500 = 2.04e-04  mcm3m1l1_cc_w_0_140_s_3_500 = 8.50e-14  mcm3m1l1_cf_w_0_140_s_3_500 = 7.11e-11
+ mcm3m1l1_ca_w_1_120_s_0_140 = 2.04e-04  mcm3m1l1_cc_w_1_120_s_0_140 = 1.10e-10  mcm3m1l1_cf_w_1_120_s_0_140 = 1.14e-11
+ mcm3m1l1_ca_w_1_120_s_0_175 = 2.04e-04  mcm3m1l1_cc_w_1_120_s_0_175 = 1.04e-10  mcm3m1l1_cf_w_1_120_s_0_175 = 1.49e-11
+ mcm3m1l1_ca_w_1_120_s_0_210 = 2.04e-04  mcm3m1l1_cc_w_1_120_s_0_210 = 9.62e-11  mcm3m1l1_cf_w_1_120_s_0_210 = 1.82e-11
+ mcm3m1l1_ca_w_1_120_s_0_280 = 2.04e-04  mcm3m1l1_cc_w_1_120_s_0_280 = 7.87e-11  mcm3m1l1_cf_w_1_120_s_0_280 = 2.44e-11
+ mcm3m1l1_ca_w_1_120_s_0_350 = 2.04e-04  mcm3m1l1_cc_w_1_120_s_0_350 = 6.33e-11  mcm3m1l1_cf_w_1_120_s_0_350 = 3.01e-11
+ mcm3m1l1_ca_w_1_120_s_0_420 = 2.04e-04  mcm3m1l1_cc_w_1_120_s_0_420 = 5.10e-11  mcm3m1l1_cf_w_1_120_s_0_420 = 3.53e-11
+ mcm3m1l1_ca_w_1_120_s_0_560 = 2.04e-04  mcm3m1l1_cc_w_1_120_s_0_560 = 3.39e-11  mcm3m1l1_cf_w_1_120_s_0_560 = 4.40e-11
+ mcm3m1l1_ca_w_1_120_s_0_840 = 2.04e-04  mcm3m1l1_cc_w_1_120_s_0_840 = 1.67e-11  mcm3m1l1_cf_w_1_120_s_0_840 = 5.61e-11
+ mcm3m1l1_ca_w_1_120_s_1_540 = 2.04e-04  mcm3m1l1_cc_w_1_120_s_1_540 = 3.40e-12  mcm3m1l1_cf_w_1_120_s_1_540 = 6.84e-11
+ mcm3m1l1_ca_w_1_120_s_3_500 = 2.04e-04  mcm3m1l1_cc_w_1_120_s_3_500 = 9.00e-14  mcm3m1l1_cf_w_1_120_s_3_500 = 7.24e-11
+ mcm4m1f_ca_w_0_140_s_0_140 = 4.91e-05  mcm4m1f_cc_w_0_140_s_0_140 = 1.20e-10  mcm4m1f_cf_w_0_140_s_0_140 = 2.88e-12
+ mcm4m1f_ca_w_0_140_s_0_175 = 4.91e-05  mcm4m1f_cc_w_0_140_s_0_175 = 1.15e-10  mcm4m1f_cf_w_0_140_s_0_175 = 3.73e-12
+ mcm4m1f_ca_w_0_140_s_0_210 = 4.91e-05  mcm4m1f_cc_w_0_140_s_0_210 = 1.09e-10  mcm4m1f_cf_w_0_140_s_0_210 = 4.59e-12
+ mcm4m1f_ca_w_0_140_s_0_280 = 4.91e-05  mcm4m1f_cc_w_0_140_s_0_280 = 9.33e-11  mcm4m1f_cf_w_0_140_s_0_280 = 6.25e-12
+ mcm4m1f_ca_w_0_140_s_0_350 = 4.91e-05  mcm4m1f_cc_w_0_140_s_0_350 = 7.98e-11  mcm4m1f_cf_w_0_140_s_0_350 = 7.88e-12
+ mcm4m1f_ca_w_0_140_s_0_420 = 4.91e-05  mcm4m1f_cc_w_0_140_s_0_420 = 6.80e-11  mcm4m1f_cf_w_0_140_s_0_420 = 9.54e-12
+ mcm4m1f_ca_w_0_140_s_0_560 = 4.91e-05  mcm4m1f_cc_w_0_140_s_0_560 = 5.23e-11  mcm4m1f_cf_w_0_140_s_0_560 = 1.26e-11
+ mcm4m1f_ca_w_0_140_s_0_840 = 4.91e-05  mcm4m1f_cc_w_0_140_s_0_840 = 3.51e-11  mcm4m1f_cf_w_0_140_s_0_840 = 1.81e-11
+ mcm4m1f_ca_w_0_140_s_1_540 = 4.91e-05  mcm4m1f_cc_w_0_140_s_1_540 = 1.62e-11  mcm4m1f_cf_w_0_140_s_1_540 = 2.85e-11
+ mcm4m1f_ca_w_0_140_s_3_500 = 4.91e-05  mcm4m1f_cc_w_0_140_s_3_500 = 2.56e-12  mcm4m1f_cf_w_0_140_s_3_500 = 3.98e-11
+ mcm4m1f_ca_w_1_120_s_0_140 = 4.91e-05  mcm4m1f_cc_w_1_120_s_0_140 = 1.37e-10  mcm4m1f_cf_w_1_120_s_0_140 = 2.94e-12
+ mcm4m1f_ca_w_1_120_s_0_175 = 4.91e-05  mcm4m1f_cc_w_1_120_s_0_175 = 1.32e-10  mcm4m1f_cf_w_1_120_s_0_175 = 3.80e-12
+ mcm4m1f_ca_w_1_120_s_0_210 = 4.91e-05  mcm4m1f_cc_w_1_120_s_0_210 = 1.24e-10  mcm4m1f_cf_w_1_120_s_0_210 = 4.64e-12
+ mcm4m1f_ca_w_1_120_s_0_280 = 4.91e-05  mcm4m1f_cc_w_1_120_s_0_280 = 1.06e-10  mcm4m1f_cf_w_1_120_s_0_280 = 6.31e-12
+ mcm4m1f_ca_w_1_120_s_0_350 = 4.91e-05  mcm4m1f_cc_w_1_120_s_0_350 = 9.02e-11  mcm4m1f_cf_w_1_120_s_0_350 = 7.95e-12
+ mcm4m1f_ca_w_1_120_s_0_420 = 4.91e-05  mcm4m1f_cc_w_1_120_s_0_420 = 7.79e-11  mcm4m1f_cf_w_1_120_s_0_420 = 9.56e-12
+ mcm4m1f_ca_w_1_120_s_0_560 = 4.91e-05  mcm4m1f_cc_w_1_120_s_0_560 = 6.02e-11  mcm4m1f_cf_w_1_120_s_0_560 = 1.27e-11
+ mcm4m1f_ca_w_1_120_s_0_840 = 4.91e-05  mcm4m1f_cc_w_1_120_s_0_840 = 4.03e-11  mcm4m1f_cf_w_1_120_s_0_840 = 1.83e-11
+ mcm4m1f_ca_w_1_120_s_1_540 = 4.91e-05  mcm4m1f_cc_w_1_120_s_1_540 = 1.87e-11  mcm4m1f_cf_w_1_120_s_1_540 = 2.94e-11
+ mcm4m1f_ca_w_1_120_s_3_500 = 4.91e-05  mcm4m1f_cc_w_1_120_s_3_500 = 3.03e-12  mcm4m1f_cf_w_1_120_s_3_500 = 4.20e-11
+ mcm4m1d_ca_w_0_140_s_0_140 = 5.81e-05  mcm4m1d_cc_w_0_140_s_0_140 = 1.17e-10  mcm4m1d_cf_w_0_140_s_0_140 = 3.40e-12
+ mcm4m1d_ca_w_0_140_s_0_175 = 5.81e-05  mcm4m1d_cc_w_0_140_s_0_175 = 1.14e-10  mcm4m1d_cf_w_0_140_s_0_175 = 4.40e-12
+ mcm4m1d_ca_w_0_140_s_0_210 = 5.81e-05  mcm4m1d_cc_w_0_140_s_0_210 = 1.07e-10  mcm4m1d_cf_w_0_140_s_0_210 = 5.41e-12
+ mcm4m1d_ca_w_0_140_s_0_280 = 5.81e-05  mcm4m1d_cc_w_0_140_s_0_280 = 9.24e-11  mcm4m1d_cf_w_0_140_s_0_280 = 7.37e-12
+ mcm4m1d_ca_w_0_140_s_0_350 = 5.81e-05  mcm4m1d_cc_w_0_140_s_0_350 = 7.83e-11  mcm4m1d_cf_w_0_140_s_0_350 = 9.29e-12
+ mcm4m1d_ca_w_0_140_s_0_420 = 5.81e-05  mcm4m1d_cc_w_0_140_s_0_420 = 6.63e-11  mcm4m1d_cf_w_0_140_s_0_420 = 1.12e-11
+ mcm4m1d_ca_w_0_140_s_0_560 = 5.81e-05  mcm4m1d_cc_w_0_140_s_0_560 = 5.04e-11  mcm4m1d_cf_w_0_140_s_0_560 = 1.47e-11
+ mcm4m1d_ca_w_0_140_s_0_840 = 5.81e-05  mcm4m1d_cc_w_0_140_s_0_840 = 3.30e-11  mcm4m1d_cf_w_0_140_s_0_840 = 2.10e-11
+ mcm4m1d_ca_w_0_140_s_1_540 = 5.81e-05  mcm4m1d_cc_w_0_140_s_1_540 = 1.42e-11  mcm4m1d_cf_w_0_140_s_1_540 = 3.22e-11
+ mcm4m1d_ca_w_0_140_s_3_500 = 5.81e-05  mcm4m1d_cc_w_0_140_s_3_500 = 1.92e-12  mcm4m1d_cf_w_0_140_s_3_500 = 4.28e-11
+ mcm4m1d_ca_w_1_120_s_0_140 = 5.81e-05  mcm4m1d_cc_w_1_120_s_0_140 = 1.35e-10  mcm4m1d_cf_w_1_120_s_0_140 = 3.50e-12
+ mcm4m1d_ca_w_1_120_s_0_175 = 5.81e-05  mcm4m1d_cc_w_1_120_s_0_175 = 1.29e-10  mcm4m1d_cf_w_1_120_s_0_175 = 4.51e-12
+ mcm4m1d_ca_w_1_120_s_0_210 = 5.81e-05  mcm4m1d_cc_w_1_120_s_0_210 = 1.22e-10  mcm4m1d_cf_w_1_120_s_0_210 = 5.51e-12
+ mcm4m1d_ca_w_1_120_s_0_280 = 5.81e-05  mcm4m1d_cc_w_1_120_s_0_280 = 1.03e-10  mcm4m1d_cf_w_1_120_s_0_280 = 7.45e-12
+ mcm4m1d_ca_w_1_120_s_0_350 = 5.81e-05  mcm4m1d_cc_w_1_120_s_0_350 = 8.73e-11  mcm4m1d_cf_w_1_120_s_0_350 = 9.38e-12
+ mcm4m1d_ca_w_1_120_s_0_420 = 5.81e-05  mcm4m1d_cc_w_1_120_s_0_420 = 7.53e-11  mcm4m1d_cf_w_1_120_s_0_420 = 1.13e-11
+ mcm4m1d_ca_w_1_120_s_0_560 = 5.81e-05  mcm4m1d_cc_w_1_120_s_0_560 = 5.72e-11  mcm4m1d_cf_w_1_120_s_0_560 = 1.49e-11
+ mcm4m1d_ca_w_1_120_s_0_840 = 5.81e-05  mcm4m1d_cc_w_1_120_s_0_840 = 3.76e-11  mcm4m1d_cf_w_1_120_s_0_840 = 2.13e-11
+ mcm4m1d_ca_w_1_120_s_1_540 = 5.81e-05  mcm4m1d_cc_w_1_120_s_1_540 = 1.65e-11  mcm4m1d_cf_w_1_120_s_1_540 = 3.31e-11
+ mcm4m1d_ca_w_1_120_s_3_500 = 5.81e-05  mcm4m1d_cc_w_1_120_s_3_500 = 2.29e-12  mcm4m1d_cf_w_1_120_s_3_500 = 4.51e-11
+ mcm4m1p1_ca_w_0_140_s_0_140 = 7.81e-05  mcm4m1p1_cc_w_0_140_s_0_140 = 1.15e-10  mcm4m1p1_cf_w_0_140_s_0_140 = 4.57e-12
+ mcm4m1p1_ca_w_0_140_s_0_175 = 7.81e-05  mcm4m1p1_cc_w_0_140_s_0_175 = 1.12e-10  mcm4m1p1_cf_w_0_140_s_0_175 = 5.92e-12
+ mcm4m1p1_ca_w_0_140_s_0_210 = 7.81e-05  mcm4m1p1_cc_w_0_140_s_0_210 = 1.05e-10  mcm4m1p1_cf_w_0_140_s_0_210 = 7.27e-12
+ mcm4m1p1_ca_w_0_140_s_0_280 = 7.81e-05  mcm4m1p1_cc_w_0_140_s_0_280 = 8.95e-11  mcm4m1p1_cf_w_0_140_s_0_280 = 9.87e-12
+ mcm4m1p1_ca_w_0_140_s_0_350 = 7.81e-05  mcm4m1p1_cc_w_0_140_s_0_350 = 7.47e-11  mcm4m1p1_cf_w_0_140_s_0_350 = 1.24e-11
+ mcm4m1p1_ca_w_0_140_s_0_420 = 7.81e-05  mcm4m1p1_cc_w_0_140_s_0_420 = 6.32e-11  mcm4m1p1_cf_w_0_140_s_0_420 = 1.49e-11
+ mcm4m1p1_ca_w_0_140_s_0_560 = 7.81e-05  mcm4m1p1_cc_w_0_140_s_0_560 = 4.68e-11  mcm4m1p1_cf_w_0_140_s_0_560 = 1.94e-11
+ mcm4m1p1_ca_w_0_140_s_0_840 = 7.81e-05  mcm4m1p1_cc_w_0_140_s_0_840 = 2.92e-11  mcm4m1p1_cf_w_0_140_s_0_840 = 2.70e-11
+ mcm4m1p1_ca_w_0_140_s_1_540 = 7.81e-05  mcm4m1p1_cc_w_0_140_s_1_540 = 1.13e-11  mcm4m1p1_cf_w_0_140_s_1_540 = 3.93e-11
+ mcm4m1p1_ca_w_0_140_s_3_500 = 7.81e-05  mcm4m1p1_cc_w_0_140_s_3_500 = 1.19e-12  mcm4m1p1_cf_w_0_140_s_3_500 = 4.85e-11
+ mcm4m1p1_ca_w_1_120_s_0_140 = 7.81e-05  mcm4m1p1_cc_w_1_120_s_0_140 = 1.30e-10  mcm4m1p1_cf_w_1_120_s_0_140 = 4.80e-12
+ mcm4m1p1_ca_w_1_120_s_0_175 = 7.81e-05  mcm4m1p1_cc_w_1_120_s_0_175 = 1.24e-10  mcm4m1p1_cf_w_1_120_s_0_175 = 6.14e-12
+ mcm4m1p1_ca_w_1_120_s_0_210 = 7.81e-05  mcm4m1p1_cc_w_1_120_s_0_210 = 1.16e-10  mcm4m1p1_cf_w_1_120_s_0_210 = 7.46e-12
+ mcm4m1p1_ca_w_1_120_s_0_280 = 7.81e-05  mcm4m1p1_cc_w_1_120_s_0_280 = 9.82e-11  mcm4m1p1_cf_w_1_120_s_0_280 = 1.01e-11
+ mcm4m1p1_ca_w_1_120_s_0_350 = 7.81e-05  mcm4m1p1_cc_w_1_120_s_0_350 = 8.29e-11  mcm4m1p1_cf_w_1_120_s_0_350 = 1.26e-11
+ mcm4m1p1_ca_w_1_120_s_0_420 = 7.81e-05  mcm4m1p1_cc_w_1_120_s_0_420 = 6.99e-11  mcm4m1p1_cf_w_1_120_s_0_420 = 1.50e-11
+ mcm4m1p1_ca_w_1_120_s_0_560 = 7.81e-05  mcm4m1p1_cc_w_1_120_s_0_560 = 5.25e-11  mcm4m1p1_cf_w_1_120_s_0_560 = 1.96e-11
+ mcm4m1p1_ca_w_1_120_s_0_840 = 7.81e-05  mcm4m1p1_cc_w_1_120_s_0_840 = 3.31e-11  mcm4m1p1_cf_w_1_120_s_0_840 = 2.74e-11
+ mcm4m1p1_ca_w_1_120_s_1_540 = 7.81e-05  mcm4m1p1_cc_w_1_120_s_1_540 = 1.32e-11  mcm4m1p1_cf_w_1_120_s_1_540 = 4.04e-11
+ mcm4m1p1_ca_w_1_120_s_3_500 = 7.81e-05  mcm4m1p1_cc_w_1_120_s_3_500 = 1.50e-12  mcm4m1p1_cf_w_1_120_s_3_500 = 5.10e-11
+ mcm4m1l1_ca_w_0_140_s_0_140 = 1.80e-04  mcm4m1l1_cc_w_0_140_s_0_140 = 1.08e-10  mcm4m1l1_cf_w_0_140_s_0_140 = 9.91e-12
+ mcm4m1l1_ca_w_0_140_s_0_175 = 1.80e-04  mcm4m1l1_cc_w_0_140_s_0_175 = 1.03e-10  mcm4m1l1_cf_w_0_140_s_0_175 = 1.30e-11
+ mcm4m1l1_ca_w_0_140_s_0_210 = 1.80e-04  mcm4m1l1_cc_w_0_140_s_0_210 = 9.50e-11  mcm4m1l1_cf_w_0_140_s_0_210 = 1.60e-11
+ mcm4m1l1_ca_w_0_140_s_0_280 = 1.80e-04  mcm4m1l1_cc_w_0_140_s_0_280 = 7.97e-11  mcm4m1l1_cf_w_0_140_s_0_280 = 2.15e-11
+ mcm4m1l1_ca_w_0_140_s_0_350 = 1.80e-04  mcm4m1l1_cc_w_0_140_s_0_350 = 6.47e-11  mcm4m1l1_cf_w_0_140_s_0_350 = 2.65e-11
+ mcm4m1l1_ca_w_0_140_s_0_420 = 1.80e-04  mcm4m1l1_cc_w_0_140_s_0_420 = 5.30e-11  mcm4m1l1_cf_w_0_140_s_0_420 = 3.12e-11
+ mcm4m1l1_ca_w_0_140_s_0_560 = 1.80e-04  mcm4m1l1_cc_w_0_140_s_0_560 = 3.72e-11  mcm4m1l1_cf_w_0_140_s_0_560 = 3.88e-11
+ mcm4m1l1_ca_w_0_140_s_0_840 = 1.80e-04  mcm4m1l1_cc_w_0_140_s_0_840 = 2.07e-11  mcm4m1l1_cf_w_0_140_s_0_840 = 4.97e-11
+ mcm4m1l1_ca_w_0_140_s_1_540 = 1.80e-04  mcm4m1l1_cc_w_0_140_s_1_540 = 6.49e-12  mcm4m1l1_cf_w_0_140_s_1_540 = 6.21e-11
+ mcm4m1l1_ca_w_0_140_s_3_500 = 1.80e-04  mcm4m1l1_cc_w_0_140_s_3_500 = 5.75e-13  mcm4m1l1_cf_w_0_140_s_3_500 = 6.84e-11
+ mcm4m1l1_ca_w_1_120_s_0_140 = 1.80e-04  mcm4m1l1_cc_w_1_120_s_0_140 = 1.19e-10  mcm4m1l1_cf_w_1_120_s_0_140 = 1.01e-11
+ mcm4m1l1_ca_w_1_120_s_0_175 = 1.80e-04  mcm4m1l1_cc_w_1_120_s_0_175 = 1.12e-10  mcm4m1l1_cf_w_1_120_s_0_175 = 1.32e-11
+ mcm4m1l1_ca_w_1_120_s_0_210 = 1.80e-04  mcm4m1l1_cc_w_1_120_s_0_210 = 1.05e-10  mcm4m1l1_cf_w_1_120_s_0_210 = 1.62e-11
+ mcm4m1l1_ca_w_1_120_s_0_280 = 1.80e-04  mcm4m1l1_cc_w_1_120_s_0_280 = 8.71e-11  mcm4m1l1_cf_w_1_120_s_0_280 = 2.17e-11
+ mcm4m1l1_ca_w_1_120_s_0_350 = 1.80e-04  mcm4m1l1_cc_w_1_120_s_0_350 = 7.16e-11  mcm4m1l1_cf_w_1_120_s_0_350 = 2.67e-11
+ mcm4m1l1_ca_w_1_120_s_0_420 = 1.80e-04  mcm4m1l1_cc_w_1_120_s_0_420 = 5.91e-11  mcm4m1l1_cf_w_1_120_s_0_420 = 3.13e-11
+ mcm4m1l1_ca_w_1_120_s_0_560 = 1.80e-04  mcm4m1l1_cc_w_1_120_s_0_560 = 4.22e-11  mcm4m1l1_cf_w_1_120_s_0_560 = 3.89e-11
+ mcm4m1l1_ca_w_1_120_s_0_840 = 1.80e-04  mcm4m1l1_cc_w_1_120_s_0_840 = 2.44e-11  mcm4m1l1_cf_w_1_120_s_0_840 = 5.01e-11
+ mcm4m1l1_ca_w_1_120_s_1_540 = 1.80e-04  mcm4m1l1_cc_w_1_120_s_1_540 = 8.26e-12  mcm4m1l1_cf_w_1_120_s_1_540 = 6.35e-11
+ mcm4m1l1_ca_w_1_120_s_3_500 = 1.80e-04  mcm4m1l1_cc_w_1_120_s_3_500 = 7.60e-13  mcm4m1l1_cf_w_1_120_s_3_500 = 7.12e-11
+ mcm5m1f_ca_w_0_140_s_0_140 = 4.24e-05  mcm5m1f_cc_w_0_140_s_0_140 = 1.21e-10  mcm5m1f_cf_w_0_140_s_0_140 = 2.49e-12
+ mcm5m1f_ca_w_0_140_s_0_175 = 4.24e-05  mcm5m1f_cc_w_0_140_s_0_175 = 1.16e-10  mcm5m1f_cf_w_0_140_s_0_175 = 3.23e-12
+ mcm5m1f_ca_w_0_140_s_0_210 = 4.24e-05  mcm5m1f_cc_w_0_140_s_0_210 = 1.10e-10  mcm5m1f_cf_w_0_140_s_0_210 = 3.96e-12
+ mcm5m1f_ca_w_0_140_s_0_280 = 4.24e-05  mcm5m1f_cc_w_0_140_s_0_280 = 9.51e-11  mcm5m1f_cf_w_0_140_s_0_280 = 5.41e-12
+ mcm5m1f_ca_w_0_140_s_0_350 = 4.24e-05  mcm5m1f_cc_w_0_140_s_0_350 = 8.13e-11  mcm5m1f_cf_w_0_140_s_0_350 = 6.83e-12
+ mcm5m1f_ca_w_0_140_s_0_420 = 4.24e-05  mcm5m1f_cc_w_0_140_s_0_420 = 6.96e-11  mcm5m1f_cf_w_0_140_s_0_420 = 8.28e-12
+ mcm5m1f_ca_w_0_140_s_0_560 = 4.24e-05  mcm5m1f_cc_w_0_140_s_0_560 = 5.42e-11  mcm5m1f_cf_w_0_140_s_0_560 = 1.09e-11
+ mcm5m1f_ca_w_0_140_s_0_840 = 4.24e-05  mcm5m1f_cc_w_0_140_s_0_840 = 3.74e-11  mcm5m1f_cf_w_0_140_s_0_840 = 1.58e-11
+ mcm5m1f_ca_w_0_140_s_1_540 = 4.24e-05  mcm5m1f_cc_w_0_140_s_1_540 = 1.88e-11  mcm5m1f_cf_w_0_140_s_1_540 = 2.53e-11
+ mcm5m1f_ca_w_0_140_s_3_500 = 4.24e-05  mcm5m1f_cc_w_0_140_s_3_500 = 4.06e-12  mcm5m1f_cf_w_0_140_s_3_500 = 3.70e-11
+ mcm5m1f_ca_w_1_120_s_0_140 = 4.24e-05  mcm5m1f_cc_w_1_120_s_0_140 = 1.40e-10  mcm5m1f_cf_w_1_120_s_0_140 = 2.56e-12
+ mcm5m1f_ca_w_1_120_s_0_175 = 4.24e-05  mcm5m1f_cc_w_1_120_s_0_175 = 1.35e-10  mcm5m1f_cf_w_1_120_s_0_175 = 3.30e-12
+ mcm5m1f_ca_w_1_120_s_0_210 = 4.24e-05  mcm5m1f_cc_w_1_120_s_0_210 = 1.28e-10  mcm5m1f_cf_w_1_120_s_0_210 = 4.03e-12
+ mcm5m1f_ca_w_1_120_s_0_280 = 4.24e-05  mcm5m1f_cc_w_1_120_s_0_280 = 1.09e-10  mcm5m1f_cf_w_1_120_s_0_280 = 5.48e-12
+ mcm5m1f_ca_w_1_120_s_0_350 = 4.24e-05  mcm5m1f_cc_w_1_120_s_0_350 = 9.44e-11  mcm5m1f_cf_w_1_120_s_0_350 = 6.90e-12
+ mcm5m1f_ca_w_1_120_s_0_420 = 4.24e-05  mcm5m1f_cc_w_1_120_s_0_420 = 8.17e-11  mcm5m1f_cf_w_1_120_s_0_420 = 8.31e-12
+ mcm5m1f_ca_w_1_120_s_0_560 = 4.24e-05  mcm5m1f_cc_w_1_120_s_0_560 = 6.39e-11  mcm5m1f_cf_w_1_120_s_0_560 = 1.10e-11
+ mcm5m1f_ca_w_1_120_s_0_840 = 4.24e-05  mcm5m1f_cc_w_1_120_s_0_840 = 4.42e-11  mcm5m1f_cf_w_1_120_s_0_840 = 1.60e-11
+ mcm5m1f_ca_w_1_120_s_1_540 = 4.24e-05  mcm5m1f_cc_w_1_120_s_1_540 = 2.26e-11  mcm5m1f_cf_w_1_120_s_1_540 = 2.60e-11
+ mcm5m1f_ca_w_1_120_s_3_500 = 4.24e-05  mcm5m1f_cc_w_1_120_s_3_500 = 5.20e-12  mcm5m1f_cf_w_1_120_s_3_500 = 3.92e-11
+ mcm5m1d_ca_w_0_140_s_0_140 = 5.14e-05  mcm5m1d_cc_w_0_140_s_0_140 = 1.18e-10  mcm5m1d_cf_w_0_140_s_0_140 = 3.01e-12
+ mcm5m1d_ca_w_0_140_s_0_175 = 5.14e-05  mcm5m1d_cc_w_0_140_s_0_175 = 1.15e-10  mcm5m1d_cf_w_0_140_s_0_175 = 3.90e-12
+ mcm5m1d_ca_w_0_140_s_0_210 = 5.14e-05  mcm5m1d_cc_w_0_140_s_0_210 = 1.08e-10  mcm5m1d_cf_w_0_140_s_0_210 = 4.79e-12
+ mcm5m1d_ca_w_0_140_s_0_280 = 5.14e-05  mcm5m1d_cc_w_0_140_s_0_280 = 9.36e-11  mcm5m1d_cf_w_0_140_s_0_280 = 6.54e-12
+ mcm5m1d_ca_w_0_140_s_0_350 = 5.14e-05  mcm5m1d_cc_w_0_140_s_0_350 = 7.91e-11  mcm5m1d_cf_w_0_140_s_0_350 = 8.23e-12
+ mcm5m1d_ca_w_0_140_s_0_420 = 5.14e-05  mcm5m1d_cc_w_0_140_s_0_420 = 6.80e-11  mcm5m1d_cf_w_0_140_s_0_420 = 9.95e-12
+ mcm5m1d_ca_w_0_140_s_0_560 = 5.14e-05  mcm5m1d_cc_w_0_140_s_0_560 = 5.22e-11  mcm5m1d_cf_w_0_140_s_0_560 = 1.31e-11
+ mcm5m1d_ca_w_0_140_s_0_840 = 5.14e-05  mcm5m1d_cc_w_0_140_s_0_840 = 3.53e-11  mcm5m1d_cf_w_0_140_s_0_840 = 1.88e-11
+ mcm5m1d_ca_w_0_140_s_1_540 = 5.14e-05  mcm5m1d_cc_w_0_140_s_1_540 = 1.67e-11  mcm5m1d_cf_w_0_140_s_1_540 = 2.92e-11
+ mcm5m1d_ca_w_0_140_s_3_500 = 5.14e-05  mcm5m1d_cc_w_0_140_s_3_500 = 3.20e-12  mcm5m1d_cf_w_0_140_s_3_500 = 4.04e-11
+ mcm5m1d_ca_w_1_120_s_0_140 = 5.14e-05  mcm5m1d_cc_w_1_120_s_0_140 = 1.38e-10  mcm5m1d_cf_w_1_120_s_0_140 = 3.11e-12
+ mcm5m1d_ca_w_1_120_s_0_175 = 5.14e-05  mcm5m1d_cc_w_1_120_s_0_175 = 1.32e-10  mcm5m1d_cf_w_1_120_s_0_175 = 4.01e-12
+ mcm5m1d_ca_w_1_120_s_0_210 = 5.14e-05  mcm5m1d_cc_w_1_120_s_0_210 = 1.25e-10  mcm5m1d_cf_w_1_120_s_0_210 = 4.90e-12
+ mcm5m1d_ca_w_1_120_s_0_280 = 5.14e-05  mcm5m1d_cc_w_1_120_s_0_280 = 1.07e-10  mcm5m1d_cf_w_1_120_s_0_280 = 6.62e-12
+ mcm5m1d_ca_w_1_120_s_0_350 = 5.14e-05  mcm5m1d_cc_w_1_120_s_0_350 = 9.08e-11  mcm5m1d_cf_w_1_120_s_0_350 = 8.33e-12
+ mcm5m1d_ca_w_1_120_s_0_420 = 5.14e-05  mcm5m1d_cc_w_1_120_s_0_420 = 7.85e-11  mcm5m1d_cf_w_1_120_s_0_420 = 1.00e-11
+ mcm5m1d_ca_w_1_120_s_0_560 = 5.14e-05  mcm5m1d_cc_w_1_120_s_0_560 = 6.11e-11  mcm5m1d_cf_w_1_120_s_0_560 = 1.32e-11
+ mcm5m1d_ca_w_1_120_s_0_840 = 5.14e-05  mcm5m1d_cc_w_1_120_s_0_840 = 4.15e-11  mcm5m1d_cf_w_1_120_s_0_840 = 1.90e-11
+ mcm5m1d_ca_w_1_120_s_1_540 = 5.14e-05  mcm5m1d_cc_w_1_120_s_1_540 = 2.02e-11  mcm5m1d_cf_w_1_120_s_1_540 = 3.00e-11
+ mcm5m1d_ca_w_1_120_s_3_500 = 5.14e-05  mcm5m1d_cc_w_1_120_s_3_500 = 4.22e-12  mcm5m1d_cf_w_1_120_s_3_500 = 4.29e-11
+ mcm5m1p1_ca_w_0_140_s_0_140 = 7.14e-05  mcm5m1p1_cc_w_0_140_s_0_140 = 1.16e-10  mcm5m1p1_cf_w_0_140_s_0_140 = 4.18e-12
+ mcm5m1p1_ca_w_0_140_s_0_175 = 7.14e-05  mcm5m1p1_cc_w_0_140_s_0_175 = 1.12e-10  mcm5m1p1_cf_w_0_140_s_0_175 = 5.42e-12
+ mcm5m1p1_ca_w_0_140_s_0_210 = 7.14e-05  mcm5m1p1_cc_w_0_140_s_0_210 = 1.06e-10  mcm5m1p1_cf_w_0_140_s_0_210 = 6.65e-12
+ mcm5m1p1_ca_w_0_140_s_0_280 = 7.14e-05  mcm5m1p1_cc_w_0_140_s_0_280 = 9.06e-11  mcm5m1p1_cf_w_0_140_s_0_280 = 9.05e-12
+ mcm5m1p1_ca_w_0_140_s_0_350 = 7.14e-05  mcm5m1p1_cc_w_0_140_s_0_350 = 7.61e-11  mcm5m1p1_cf_w_0_140_s_0_350 = 1.13e-11
+ mcm5m1p1_ca_w_0_140_s_0_420 = 7.14e-05  mcm5m1p1_cc_w_0_140_s_0_420 = 6.43e-11  mcm5m1p1_cf_w_0_140_s_0_420 = 1.36e-11
+ mcm5m1p1_ca_w_0_140_s_0_560 = 7.14e-05  mcm5m1p1_cc_w_0_140_s_0_560 = 4.87e-11  mcm5m1p1_cf_w_0_140_s_0_560 = 1.78e-11
+ mcm5m1p1_ca_w_0_140_s_0_840 = 7.14e-05  mcm5m1p1_cc_w_0_140_s_0_840 = 3.14e-11  mcm5m1p1_cf_w_0_140_s_0_840 = 2.48e-11
+ mcm5m1p1_ca_w_0_140_s_1_540 = 7.14e-05  mcm5m1p1_cc_w_0_140_s_1_540 = 1.35e-11  mcm5m1p1_cf_w_0_140_s_1_540 = 3.66e-11
+ mcm5m1p1_ca_w_0_140_s_3_500 = 7.14e-05  mcm5m1p1_cc_w_0_140_s_3_500 = 2.20e-12  mcm5m1p1_cf_w_0_140_s_3_500 = 4.67e-11
+ mcm5m1p1_ca_w_1_120_s_0_140 = 7.14e-05  mcm5m1p1_cc_w_1_120_s_0_140 = 1.32e-10  mcm5m1p1_cf_w_1_120_s_0_140 = 4.42e-12
+ mcm5m1p1_ca_w_1_120_s_0_175 = 7.14e-05  mcm5m1p1_cc_w_1_120_s_0_175 = 1.27e-10  mcm5m1p1_cf_w_1_120_s_0_175 = 5.65e-12
+ mcm5m1p1_ca_w_1_120_s_0_210 = 7.14e-05  mcm5m1p1_cc_w_1_120_s_0_210 = 1.20e-10  mcm5m1p1_cf_w_1_120_s_0_210 = 6.86e-12
+ mcm5m1p1_ca_w_1_120_s_0_280 = 7.14e-05  mcm5m1p1_cc_w_1_120_s_0_280 = 1.02e-10  mcm5m1p1_cf_w_1_120_s_0_280 = 9.24e-12
+ mcm5m1p1_ca_w_1_120_s_0_350 = 7.14e-05  mcm5m1p1_cc_w_1_120_s_0_350 = 8.63e-11  mcm5m1p1_cf_w_1_120_s_0_350 = 1.16e-11
+ mcm5m1p1_ca_w_1_120_s_0_420 = 7.14e-05  mcm5m1p1_cc_w_1_120_s_0_420 = 7.36e-11  mcm5m1p1_cf_w_1_120_s_0_420 = 1.38e-11
+ mcm5m1p1_ca_w_1_120_s_0_560 = 7.14e-05  mcm5m1p1_cc_w_1_120_s_0_560 = 5.62e-11  mcm5m1p1_cf_w_1_120_s_0_560 = 1.80e-11
+ mcm5m1p1_ca_w_1_120_s_0_840 = 7.14e-05  mcm5m1p1_cc_w_1_120_s_0_840 = 3.69e-11  mcm5m1p1_cf_w_1_120_s_0_840 = 2.51e-11
+ mcm5m1p1_ca_w_1_120_s_1_540 = 7.14e-05  mcm5m1p1_cc_w_1_120_s_1_540 = 1.68e-11  mcm5m1p1_cf_w_1_120_s_1_540 = 3.76e-11
+ mcm5m1p1_ca_w_1_120_s_3_500 = 7.14e-05  mcm5m1p1_cc_w_1_120_s_3_500 = 3.02e-12  mcm5m1p1_cf_w_1_120_s_3_500 = 4.96e-11
+ mcm5m1l1_ca_w_0_140_s_0_140 = 1.73e-04  mcm5m1l1_cc_w_0_140_s_0_140 = 1.09e-10  mcm5m1l1_cf_w_0_140_s_0_140 = 9.51e-12
+ mcm5m1l1_ca_w_0_140_s_0_175 = 1.73e-04  mcm5m1l1_cc_w_0_140_s_0_175 = 1.04e-10  mcm5m1l1_cf_w_0_140_s_0_175 = 1.25e-11
+ mcm5m1l1_ca_w_0_140_s_0_210 = 1.73e-04  mcm5m1l1_cc_w_0_140_s_0_210 = 9.59e-11  mcm5m1l1_cf_w_0_140_s_0_210 = 1.54e-11
+ mcm5m1l1_ca_w_0_140_s_0_280 = 1.73e-04  mcm5m1l1_cc_w_0_140_s_0_280 = 8.04e-11  mcm5m1l1_cf_w_0_140_s_0_280 = 2.07e-11
+ mcm5m1l1_ca_w_0_140_s_0_350 = 1.73e-04  mcm5m1l1_cc_w_0_140_s_0_350 = 6.61e-11  mcm5m1l1_cf_w_0_140_s_0_350 = 2.55e-11
+ mcm5m1l1_ca_w_0_140_s_0_420 = 1.73e-04  mcm5m1l1_cc_w_0_140_s_0_420 = 5.46e-11  mcm5m1l1_cf_w_0_140_s_0_420 = 3.00e-11
+ mcm5m1l1_ca_w_0_140_s_0_560 = 1.73e-04  mcm5m1l1_cc_w_0_140_s_0_560 = 3.89e-11  mcm5m1l1_cf_w_0_140_s_0_560 = 3.72e-11
+ mcm5m1l1_ca_w_0_140_s_0_840 = 1.73e-04  mcm5m1l1_cc_w_0_140_s_0_840 = 2.28e-11  mcm5m1l1_cf_w_0_140_s_0_840 = 4.77e-11
+ mcm5m1l1_ca_w_0_140_s_1_540 = 1.73e-04  mcm5m1l1_cc_w_0_140_s_1_540 = 8.19e-12  mcm5m1l1_cf_w_0_140_s_1_540 = 6.02e-11
+ mcm5m1l1_ca_w_0_140_s_3_500 = 1.73e-04  mcm5m1l1_cc_w_0_140_s_3_500 = 1.05e-12  mcm5m1l1_cf_w_0_140_s_3_500 = 6.75e-11
+ mcm5m1l1_ca_w_1_120_s_0_140 = 1.73e-04  mcm5m1l1_cc_w_1_120_s_0_140 = 1.22e-10  mcm5m1l1_cf_w_1_120_s_0_140 = 9.73e-12
+ mcm5m1l1_ca_w_1_120_s_0_175 = 1.73e-04  mcm5m1l1_cc_w_1_120_s_0_175 = 1.15e-10  mcm5m1l1_cf_w_1_120_s_0_175 = 1.27e-11
+ mcm5m1l1_ca_w_1_120_s_0_210 = 1.73e-04  mcm5m1l1_cc_w_1_120_s_0_210 = 1.08e-10  mcm5m1l1_cf_w_1_120_s_0_210 = 1.56e-11
+ mcm5m1l1_ca_w_1_120_s_0_280 = 1.73e-04  mcm5m1l1_cc_w_1_120_s_0_280 = 9.04e-11  mcm5m1l1_cf_w_1_120_s_0_280 = 2.09e-11
+ mcm5m1l1_ca_w_1_120_s_0_350 = 1.73e-04  mcm5m1l1_cc_w_1_120_s_0_350 = 7.49e-11  mcm5m1l1_cf_w_1_120_s_0_350 = 2.57e-11
+ mcm5m1l1_ca_w_1_120_s_0_420 = 1.73e-04  mcm5m1l1_cc_w_1_120_s_0_420 = 6.26e-11  mcm5m1l1_cf_w_1_120_s_0_420 = 3.01e-11
+ mcm5m1l1_ca_w_1_120_s_0_560 = 1.73e-04  mcm5m1l1_cc_w_1_120_s_0_560 = 4.58e-11  mcm5m1l1_cf_w_1_120_s_0_560 = 3.74e-11
+ mcm5m1l1_ca_w_1_120_s_0_840 = 1.73e-04  mcm5m1l1_cc_w_1_120_s_0_840 = 2.81e-11  mcm5m1l1_cf_w_1_120_s_0_840 = 4.81e-11
+ mcm5m1l1_ca_w_1_120_s_1_540 = 1.73e-04  mcm5m1l1_cc_w_1_120_s_1_540 = 1.13e-11  mcm5m1l1_cf_w_1_120_s_1_540 = 6.16e-11
+ mcm5m1l1_ca_w_1_120_s_3_500 = 1.73e-04  mcm5m1l1_cc_w_1_120_s_3_500 = 1.73e-12  mcm5m1l1_cf_w_1_120_s_3_500 = 7.11e-11
+ mcrdlm1f_ca_w_0_140_s_0_140 = 3.56e-05  mcrdlm1f_cc_w_0_140_s_0_140 = 1.21e-10  mcrdlm1f_cf_w_0_140_s_0_140 = 2.09e-12
+ mcrdlm1f_ca_w_0_140_s_0_175 = 3.56e-05  mcrdlm1f_cc_w_0_140_s_0_175 = 1.16e-10  mcrdlm1f_cf_w_0_140_s_0_175 = 2.71e-12
+ mcrdlm1f_ca_w_0_140_s_0_210 = 3.56e-05  mcrdlm1f_cc_w_0_140_s_0_210 = 1.11e-10  mcrdlm1f_cf_w_0_140_s_0_210 = 3.33e-12
+ mcrdlm1f_ca_w_0_140_s_0_280 = 3.56e-05  mcrdlm1f_cc_w_0_140_s_0_280 = 9.51e-11  mcrdlm1f_cf_w_0_140_s_0_280 = 4.54e-12
+ mcrdlm1f_ca_w_0_140_s_0_350 = 3.56e-05  mcrdlm1f_cc_w_0_140_s_0_350 = 8.19e-11  mcrdlm1f_cf_w_0_140_s_0_350 = 5.73e-12
+ mcrdlm1f_ca_w_0_140_s_0_420 = 3.56e-05  mcrdlm1f_cc_w_0_140_s_0_420 = 7.10e-11  mcrdlm1f_cf_w_0_140_s_0_420 = 6.95e-12
+ mcrdlm1f_ca_w_0_140_s_0_560 = 3.56e-05  mcrdlm1f_cc_w_0_140_s_0_560 = 5.63e-11  mcrdlm1f_cf_w_0_140_s_0_560 = 9.19e-12
+ mcrdlm1f_ca_w_0_140_s_0_840 = 3.56e-05  mcrdlm1f_cc_w_0_140_s_0_840 = 4.00e-11  mcrdlm1f_cf_w_0_140_s_0_840 = 1.33e-11
+ mcrdlm1f_ca_w_0_140_s_1_540 = 3.56e-05  mcrdlm1f_cc_w_0_140_s_1_540 = 2.21e-11  mcrdlm1f_cf_w_0_140_s_1_540 = 2.17e-11
+ mcrdlm1f_ca_w_0_140_s_3_500 = 3.56e-05  mcrdlm1f_cc_w_0_140_s_3_500 = 6.92e-12  mcrdlm1f_cf_w_0_140_s_3_500 = 3.33e-11
+ mcrdlm1f_ca_w_1_120_s_0_140 = 3.56e-05  mcrdlm1f_cc_w_1_120_s_0_140 = 1.44e-10  mcrdlm1f_cf_w_1_120_s_0_140 = 2.16e-12
+ mcrdlm1f_ca_w_1_120_s_0_175 = 3.56e-05  mcrdlm1f_cc_w_1_120_s_0_175 = 1.37e-10  mcrdlm1f_cf_w_1_120_s_0_175 = 2.78e-12
+ mcrdlm1f_ca_w_1_120_s_0_210 = 3.56e-05  mcrdlm1f_cc_w_1_120_s_0_210 = 1.30e-10  mcrdlm1f_cf_w_1_120_s_0_210 = 3.40e-12
+ mcrdlm1f_ca_w_1_120_s_0_280 = 3.56e-05  mcrdlm1f_cc_w_1_120_s_0_280 = 1.13e-10  mcrdlm1f_cf_w_1_120_s_0_280 = 4.61e-12
+ mcrdlm1f_ca_w_1_120_s_0_350 = 3.56e-05  mcrdlm1f_cc_w_1_120_s_0_350 = 9.77e-11  mcrdlm1f_cf_w_1_120_s_0_350 = 5.81e-12
+ mcrdlm1f_ca_w_1_120_s_0_420 = 3.56e-05  mcrdlm1f_cc_w_1_120_s_0_420 = 8.55e-11  mcrdlm1f_cf_w_1_120_s_0_420 = 6.99e-12
+ mcrdlm1f_ca_w_1_120_s_0_560 = 3.56e-05  mcrdlm1f_cc_w_1_120_s_0_560 = 6.82e-11  mcrdlm1f_cf_w_1_120_s_0_560 = 9.24e-12
+ mcrdlm1f_ca_w_1_120_s_0_840 = 3.56e-05  mcrdlm1f_cc_w_1_120_s_0_840 = 4.93e-11  mcrdlm1f_cf_w_1_120_s_0_840 = 1.35e-11
+ mcrdlm1f_ca_w_1_120_s_1_540 = 3.56e-05  mcrdlm1f_cc_w_1_120_s_1_540 = 2.83e-11  mcrdlm1f_cf_w_1_120_s_1_540 = 2.22e-11
+ mcrdlm1f_ca_w_1_120_s_3_500 = 3.56e-05  mcrdlm1f_cc_w_1_120_s_3_500 = 9.73e-12  mcrdlm1f_cf_w_1_120_s_3_500 = 3.55e-11
+ mcrdlm1d_ca_w_0_140_s_0_140 = 4.45e-05  mcrdlm1d_cc_w_0_140_s_0_140 = 1.19e-10  mcrdlm1d_cf_w_0_140_s_0_140 = 2.61e-12
+ mcrdlm1d_ca_w_0_140_s_0_175 = 4.45e-05  mcrdlm1d_cc_w_0_140_s_0_175 = 1.16e-10  mcrdlm1d_cf_w_0_140_s_0_175 = 3.38e-12
+ mcrdlm1d_ca_w_0_140_s_0_210 = 4.45e-05  mcrdlm1d_cc_w_0_140_s_0_210 = 1.10e-10  mcrdlm1d_cf_w_0_140_s_0_210 = 4.16e-12
+ mcrdlm1d_ca_w_0_140_s_0_280 = 4.45e-05  mcrdlm1d_cc_w_0_140_s_0_280 = 9.38e-11  mcrdlm1d_cf_w_0_140_s_0_280 = 5.67e-12
+ mcrdlm1d_ca_w_0_140_s_0_350 = 4.45e-05  mcrdlm1d_cc_w_0_140_s_0_350 = 8.04e-11  mcrdlm1d_cf_w_0_140_s_0_350 = 7.14e-12
+ mcrdlm1d_ca_w_0_140_s_0_420 = 4.45e-05  mcrdlm1d_cc_w_0_140_s_0_420 = 6.94e-11  mcrdlm1d_cf_w_0_140_s_0_420 = 8.62e-12
+ mcrdlm1d_ca_w_0_140_s_0_560 = 4.45e-05  mcrdlm1d_cc_w_0_140_s_0_560 = 5.42e-11  mcrdlm1d_cf_w_0_140_s_0_560 = 1.13e-11
+ mcrdlm1d_ca_w_0_140_s_0_840 = 4.45e-05  mcrdlm1d_cc_w_0_140_s_0_840 = 3.78e-11  mcrdlm1d_cf_w_0_140_s_0_840 = 1.63e-11
+ mcrdlm1d_ca_w_0_140_s_1_540 = 4.45e-05  mcrdlm1d_cc_w_0_140_s_1_540 = 1.99e-11  mcrdlm1d_cf_w_0_140_s_1_540 = 2.57e-11
+ mcrdlm1d_ca_w_0_140_s_3_500 = 4.45e-05  mcrdlm1d_cc_w_0_140_s_3_500 = 5.64e-12  mcrdlm1d_cf_w_0_140_s_3_500 = 3.72e-11
+ mcrdlm1d_ca_w_1_120_s_0_140 = 4.45e-05  mcrdlm1d_cc_w_1_120_s_0_140 = 1.41e-10  mcrdlm1d_cf_w_1_120_s_0_140 = 2.72e-12
+ mcrdlm1d_ca_w_1_120_s_0_175 = 4.45e-05  mcrdlm1d_cc_w_1_120_s_0_175 = 1.35e-10  mcrdlm1d_cf_w_1_120_s_0_175 = 3.48e-12
+ mcrdlm1d_ca_w_1_120_s_0_210 = 4.45e-05  mcrdlm1d_cc_w_1_120_s_0_210 = 1.27e-10  mcrdlm1d_cf_w_1_120_s_0_210 = 4.25e-12
+ mcrdlm1d_ca_w_1_120_s_0_280 = 4.45e-05  mcrdlm1d_cc_w_1_120_s_0_280 = 1.10e-10  mcrdlm1d_cf_w_1_120_s_0_280 = 5.76e-12
+ mcrdlm1d_ca_w_1_120_s_0_350 = 4.45e-05  mcrdlm1d_cc_w_1_120_s_0_350 = 9.53e-11  mcrdlm1d_cf_w_1_120_s_0_350 = 7.23e-12
+ mcrdlm1d_ca_w_1_120_s_0_420 = 4.45e-05  mcrdlm1d_cc_w_1_120_s_0_420 = 8.30e-11  mcrdlm1d_cf_w_1_120_s_0_420 = 8.68e-12
+ mcrdlm1d_ca_w_1_120_s_0_560 = 4.45e-05  mcrdlm1d_cc_w_1_120_s_0_560 = 6.53e-11  mcrdlm1d_cf_w_1_120_s_0_560 = 1.14e-11
+ mcrdlm1d_ca_w_1_120_s_0_840 = 4.45e-05  mcrdlm1d_cc_w_1_120_s_0_840 = 4.64e-11  mcrdlm1d_cf_w_1_120_s_0_840 = 1.65e-11
+ mcrdlm1d_ca_w_1_120_s_1_540 = 4.45e-05  mcrdlm1d_cc_w_1_120_s_1_540 = 2.57e-11  mcrdlm1d_cf_w_1_120_s_1_540 = 2.64e-11
+ mcrdlm1d_ca_w_1_120_s_3_500 = 4.45e-05  mcrdlm1d_cc_w_1_120_s_3_500 = 8.31e-12  mcrdlm1d_cf_w_1_120_s_3_500 = 3.98e-11
+ mcrdlm1p1_ca_w_0_140_s_0_140 = 6.45e-05  mcrdlm1p1_cc_w_0_140_s_0_140 = 1.17e-10  mcrdlm1p1_cf_w_0_140_s_0_140 = 3.77e-12
+ mcrdlm1p1_ca_w_0_140_s_0_175 = 6.45e-05  mcrdlm1p1_cc_w_0_140_s_0_175 = 1.13e-10  mcrdlm1p1_cf_w_0_140_s_0_175 = 4.89e-12
+ mcrdlm1p1_ca_w_0_140_s_0_210 = 6.45e-05  mcrdlm1p1_cc_w_0_140_s_0_210 = 1.07e-10  mcrdlm1p1_cf_w_0_140_s_0_210 = 6.02e-12
+ mcrdlm1p1_ca_w_0_140_s_0_280 = 6.45e-05  mcrdlm1p1_cc_w_0_140_s_0_280 = 9.08e-11  mcrdlm1p1_cf_w_0_140_s_0_280 = 8.17e-12
+ mcrdlm1p1_ca_w_0_140_s_0_350 = 6.45e-05  mcrdlm1p1_cc_w_0_140_s_0_350 = 7.74e-11  mcrdlm1p1_cf_w_0_140_s_0_350 = 1.02e-11
+ mcrdlm1p1_ca_w_0_140_s_0_420 = 6.45e-05  mcrdlm1p1_cc_w_0_140_s_0_420 = 6.57e-11  mcrdlm1p1_cf_w_0_140_s_0_420 = 1.23e-11
+ mcrdlm1p1_ca_w_0_140_s_0_560 = 6.45e-05  mcrdlm1p1_cc_w_0_140_s_0_560 = 5.04e-11  mcrdlm1p1_cf_w_0_140_s_0_560 = 1.60e-11
+ mcrdlm1p1_ca_w_0_140_s_0_840 = 6.45e-05  mcrdlm1p1_cc_w_0_140_s_0_840 = 3.38e-11  mcrdlm1p1_cf_w_0_140_s_0_840 = 2.25e-11
+ mcrdlm1p1_ca_w_0_140_s_1_540 = 6.45e-05  mcrdlm1p1_cc_w_0_140_s_1_540 = 1.65e-11  mcrdlm1p1_cf_w_0_140_s_1_540 = 3.35e-11
+ mcrdlm1p1_ca_w_0_140_s_3_500 = 6.45e-05  mcrdlm1p1_cc_w_0_140_s_3_500 = 4.13e-12  mcrdlm1p1_cf_w_0_140_s_3_500 = 4.43e-11
+ mcrdlm1p1_ca_w_1_120_s_0_140 = 6.45e-05  mcrdlm1p1_cc_w_1_120_s_0_140 = 1.36e-10  mcrdlm1p1_cf_w_1_120_s_0_140 = 3.99e-12
+ mcrdlm1p1_ca_w_1_120_s_0_175 = 6.45e-05  mcrdlm1p1_cc_w_1_120_s_0_175 = 1.30e-10  mcrdlm1p1_cf_w_1_120_s_0_175 = 5.12e-12
+ mcrdlm1p1_ca_w_1_120_s_0_210 = 6.45e-05  mcrdlm1p1_cc_w_1_120_s_0_210 = 1.23e-10  mcrdlm1p1_cf_w_1_120_s_0_210 = 6.23e-12
+ mcrdlm1p1_ca_w_1_120_s_0_280 = 6.45e-05  mcrdlm1p1_cc_w_1_120_s_0_280 = 1.05e-10  mcrdlm1p1_cf_w_1_120_s_0_280 = 8.37e-12
+ mcrdlm1p1_ca_w_1_120_s_0_350 = 6.45e-05  mcrdlm1p1_cc_w_1_120_s_0_350 = 9.04e-11  mcrdlm1p1_cf_w_1_120_s_0_350 = 1.05e-11
+ mcrdlm1p1_ca_w_1_120_s_0_420 = 6.45e-05  mcrdlm1p1_cc_w_1_120_s_0_420 = 7.80e-11  mcrdlm1p1_cf_w_1_120_s_0_420 = 1.25e-11
+ mcrdlm1p1_ca_w_1_120_s_0_560 = 6.45e-05  mcrdlm1p1_cc_w_1_120_s_0_560 = 6.07e-11  mcrdlm1p1_cf_w_1_120_s_0_560 = 1.62e-11
+ mcrdlm1p1_ca_w_1_120_s_0_840 = 6.45e-05  mcrdlm1p1_cc_w_1_120_s_0_840 = 4.20e-11  mcrdlm1p1_cf_w_1_120_s_0_840 = 2.27e-11
+ mcrdlm1p1_ca_w_1_120_s_1_540 = 6.45e-05  mcrdlm1p1_cc_w_1_120_s_1_540 = 2.20e-11  mcrdlm1p1_cf_w_1_120_s_1_540 = 3.44e-11
+ mcrdlm1p1_ca_w_1_120_s_3_500 = 6.45e-05  mcrdlm1p1_cc_w_1_120_s_3_500 = 6.58e-12  mcrdlm1p1_cf_w_1_120_s_3_500 = 4.73e-11
+ mcrdlm1l1_ca_w_0_140_s_0_140 = 1.67e-04  mcrdlm1l1_cc_w_0_140_s_0_140 = 1.09e-10  mcrdlm1l1_cf_w_0_140_s_0_140 = 9.10e-12
+ mcrdlm1l1_ca_w_0_140_s_0_175 = 1.67e-04  mcrdlm1l1_cc_w_0_140_s_0_175 = 1.04e-10  mcrdlm1l1_cf_w_0_140_s_0_175 = 1.20e-11
+ mcrdlm1l1_ca_w_0_140_s_0_210 = 1.67e-04  mcrdlm1l1_cc_w_0_140_s_0_210 = 9.70e-11  mcrdlm1l1_cf_w_0_140_s_0_210 = 1.47e-11
+ mcrdlm1l1_ca_w_0_140_s_0_280 = 1.67e-04  mcrdlm1l1_cc_w_0_140_s_0_280 = 8.14e-11  mcrdlm1l1_cf_w_0_140_s_0_280 = 1.98e-11
+ mcrdlm1l1_ca_w_0_140_s_0_350 = 1.67e-04  mcrdlm1l1_cc_w_0_140_s_0_350 = 6.70e-11  mcrdlm1l1_cf_w_0_140_s_0_350 = 2.43e-11
+ mcrdlm1l1_ca_w_0_140_s_0_420 = 1.67e-04  mcrdlm1l1_cc_w_0_140_s_0_420 = 5.57e-11  mcrdlm1l1_cf_w_0_140_s_0_420 = 2.86e-11
+ mcrdlm1l1_ca_w_0_140_s_0_560 = 1.67e-04  mcrdlm1l1_cc_w_0_140_s_0_560 = 4.07e-11  mcrdlm1l1_cf_w_0_140_s_0_560 = 3.55e-11
+ mcrdlm1l1_ca_w_0_140_s_0_840 = 1.67e-04  mcrdlm1l1_cc_w_0_140_s_0_840 = 2.50e-11  mcrdlm1l1_cf_w_0_140_s_0_840 = 4.54e-11
+ mcrdlm1l1_ca_w_0_140_s_1_540 = 1.67e-04  mcrdlm1l1_cc_w_0_140_s_1_540 = 1.04e-11  mcrdlm1l1_cf_w_0_140_s_1_540 = 5.79e-11
+ mcrdlm1l1_ca_w_0_140_s_3_500 = 1.67e-04  mcrdlm1l1_cc_w_0_140_s_3_500 = 2.23e-12  mcrdlm1l1_cf_w_0_140_s_3_500 = 6.62e-11
+ mcrdlm1l1_ca_w_1_120_s_0_140 = 1.67e-04  mcrdlm1l1_cc_w_1_120_s_0_140 = 1.26e-10  mcrdlm1l1_cf_w_1_120_s_0_140 = 9.34e-12
+ mcrdlm1l1_ca_w_1_120_s_0_175 = 1.67e-04  mcrdlm1l1_cc_w_1_120_s_0_175 = 1.19e-10  mcrdlm1l1_cf_w_1_120_s_0_175 = 1.22e-11
+ mcrdlm1l1_ca_w_1_120_s_0_210 = 1.67e-04  mcrdlm1l1_cc_w_1_120_s_0_210 = 1.11e-10  mcrdlm1l1_cf_w_1_120_s_0_210 = 1.49e-11
+ mcrdlm1l1_ca_w_1_120_s_0_280 = 1.67e-04  mcrdlm1l1_cc_w_1_120_s_0_280 = 9.38e-11  mcrdlm1l1_cf_w_1_120_s_0_280 = 2.00e-11
+ mcrdlm1l1_ca_w_1_120_s_0_350 = 1.67e-04  mcrdlm1l1_cc_w_1_120_s_0_350 = 7.89e-11  mcrdlm1l1_cf_w_1_120_s_0_350 = 2.46e-11
+ mcrdlm1l1_ca_w_1_120_s_0_420 = 1.67e-04  mcrdlm1l1_cc_w_1_120_s_0_420 = 6.68e-11  mcrdlm1l1_cf_w_1_120_s_0_420 = 2.87e-11
+ mcrdlm1l1_ca_w_1_120_s_0_560 = 1.67e-04  mcrdlm1l1_cc_w_1_120_s_0_560 = 5.03e-11  mcrdlm1l1_cf_w_1_120_s_0_560 = 3.57e-11
+ mcrdlm1l1_ca_w_1_120_s_0_840 = 1.67e-04  mcrdlm1l1_cc_w_1_120_s_0_840 = 3.28e-11  mcrdlm1l1_cf_w_1_120_s_0_840 = 4.58e-11
+ mcrdlm1l1_ca_w_1_120_s_1_540 = 1.67e-04  mcrdlm1l1_cc_w_1_120_s_1_540 = 1.58e-11  mcrdlm1l1_cf_w_1_120_s_1_540 = 5.93e-11
+ mcrdlm1l1_ca_w_1_120_s_3_500 = 1.67e-04  mcrdlm1l1_cc_w_1_120_s_3_500 = 4.29e-12  mcrdlm1l1_cf_w_1_120_s_3_500 = 7.03e-11
+ mcm3m2f_ca_w_0_140_s_0_140 = 1.34e-04  mcm3m2f_cc_w_0_140_s_0_140 = 1.11e-10  mcm3m2f_cf_w_0_140_s_0_140 = 7.40e-12
+ mcm3m2f_ca_w_0_140_s_0_175 = 1.34e-04  mcm3m2f_cc_w_0_140_s_0_175 = 1.06e-10  mcm3m2f_cf_w_0_140_s_0_175 = 9.44e-12
+ mcm3m2f_ca_w_0_140_s_0_210 = 1.34e-04  mcm3m2f_cc_w_0_140_s_0_210 = 9.90e-11  mcm3m2f_cf_w_0_140_s_0_210 = 1.14e-11
+ mcm3m2f_ca_w_0_140_s_0_280 = 1.34e-04  mcm3m2f_cc_w_0_140_s_0_280 = 8.32e-11  mcm3m2f_cf_w_0_140_s_0_280 = 1.52e-11
+ mcm3m2f_ca_w_0_140_s_0_350 = 1.34e-04  mcm3m2f_cc_w_0_140_s_0_350 = 6.84e-11  mcm3m2f_cf_w_0_140_s_0_350 = 1.88e-11
+ mcm3m2f_ca_w_0_140_s_0_420 = 1.34e-04  mcm3m2f_cc_w_0_140_s_0_420 = 5.69e-11  mcm3m2f_cf_w_0_140_s_0_420 = 2.23e-11
+ mcm3m2f_ca_w_0_140_s_0_560 = 1.34e-04  mcm3m2f_cc_w_0_140_s_0_560 = 4.04e-11  mcm3m2f_cf_w_0_140_s_0_560 = 2.82e-11
+ mcm3m2f_ca_w_0_140_s_0_840 = 1.34e-04  mcm3m2f_cc_w_0_140_s_0_840 = 2.33e-11  mcm3m2f_cf_w_0_140_s_0_840 = 3.74e-11
+ mcm3m2f_ca_w_0_140_s_1_540 = 1.34e-04  mcm3m2f_cc_w_0_140_s_1_540 = 7.49e-12  mcm3m2f_cf_w_0_140_s_1_540 = 4.97e-11
+ mcm3m2f_ca_w_0_140_s_3_500 = 1.34e-04  mcm3m2f_cc_w_0_140_s_3_500 = 5.35e-13  mcm3m2f_cf_w_0_140_s_3_500 = 5.65e-11
+ mcm3m2f_ca_w_1_120_s_0_140 = 1.34e-04  mcm3m2f_cc_w_1_120_s_0_140 = 1.22e-10  mcm3m2f_cf_w_1_120_s_0_140 = 7.42e-12
+ mcm3m2f_ca_w_1_120_s_0_175 = 1.34e-04  mcm3m2f_cc_w_1_120_s_0_175 = 1.15e-10  mcm3m2f_cf_w_1_120_s_0_175 = 9.48e-12
+ mcm3m2f_ca_w_1_120_s_0_210 = 1.34e-04  mcm3m2f_cc_w_1_120_s_0_210 = 1.07e-10  mcm3m2f_cf_w_1_120_s_0_210 = 1.15e-11
+ mcm3m2f_ca_w_1_120_s_0_280 = 1.34e-04  mcm3m2f_cc_w_1_120_s_0_280 = 8.94e-11  mcm3m2f_cf_w_1_120_s_0_280 = 1.53e-11
+ mcm3m2f_ca_w_1_120_s_0_350 = 1.34e-04  mcm3m2f_cc_w_1_120_s_0_350 = 7.40e-11  mcm3m2f_cf_w_1_120_s_0_350 = 1.88e-11
+ mcm3m2f_ca_w_1_120_s_0_420 = 1.34e-04  mcm3m2f_cc_w_1_120_s_0_420 = 6.18e-11  mcm3m2f_cf_w_1_120_s_0_420 = 2.22e-11
+ mcm3m2f_ca_w_1_120_s_0_560 = 1.34e-04  mcm3m2f_cc_w_1_120_s_0_560 = 4.44e-11  mcm3m2f_cf_w_1_120_s_0_560 = 2.83e-11
+ mcm3m2f_ca_w_1_120_s_0_840 = 1.34e-04  mcm3m2f_cc_w_1_120_s_0_840 = 2.60e-11  mcm3m2f_cf_w_1_120_s_0_840 = 3.77e-11
+ mcm3m2f_ca_w_1_120_s_1_540 = 1.34e-04  mcm3m2f_cc_w_1_120_s_1_540 = 8.70e-12  mcm3m2f_cf_w_1_120_s_1_540 = 5.06e-11
+ mcm3m2f_ca_w_1_120_s_3_500 = 1.34e-04  mcm3m2f_cc_w_1_120_s_3_500 = 6.30e-13  mcm3m2f_cf_w_1_120_s_3_500 = 5.83e-11
+ mcm3m2d_ca_w_0_140_s_0_140 = 1.37e-04  mcm3m2d_cc_w_0_140_s_0_140 = 1.10e-10  mcm3m2d_cf_w_0_140_s_0_140 = 7.61e-12
+ mcm3m2d_ca_w_0_140_s_0_175 = 1.37e-04  mcm3m2d_cc_w_0_140_s_0_175 = 1.05e-10  mcm3m2d_cf_w_0_140_s_0_175 = 9.73e-12
+ mcm3m2d_ca_w_0_140_s_0_210 = 1.37e-04  mcm3m2d_cc_w_0_140_s_0_210 = 9.85e-11  mcm3m2d_cf_w_0_140_s_0_210 = 1.18e-11
+ mcm3m2d_ca_w_0_140_s_0_280 = 1.37e-04  mcm3m2d_cc_w_0_140_s_0_280 = 8.23e-11  mcm3m2d_cf_w_0_140_s_0_280 = 1.57e-11
+ mcm3m2d_ca_w_0_140_s_0_350 = 1.37e-04  mcm3m2d_cc_w_0_140_s_0_350 = 6.74e-11  mcm3m2d_cf_w_0_140_s_0_350 = 1.93e-11
+ mcm3m2d_ca_w_0_140_s_0_420 = 1.37e-04  mcm3m2d_cc_w_0_140_s_0_420 = 5.59e-11  mcm3m2d_cf_w_0_140_s_0_420 = 2.29e-11
+ mcm3m2d_ca_w_0_140_s_0_560 = 1.37e-04  mcm3m2d_cc_w_0_140_s_0_560 = 3.95e-11  mcm3m2d_cf_w_0_140_s_0_560 = 2.91e-11
+ mcm3m2d_ca_w_0_140_s_0_840 = 1.37e-04  mcm3m2d_cc_w_0_140_s_0_840 = 2.23e-11  mcm3m2d_cf_w_0_140_s_0_840 = 3.86e-11
+ mcm3m2d_ca_w_0_140_s_1_540 = 1.37e-04  mcm3m2d_cc_w_0_140_s_1_540 = 6.65e-12  mcm3m2d_cf_w_0_140_s_1_540 = 5.09e-11
+ mcm3m2d_ca_w_0_140_s_3_500 = 1.37e-04  mcm3m2d_cc_w_0_140_s_3_500 = 4.10e-13  mcm3m2d_cf_w_0_140_s_3_500 = 5.70e-11
+ mcm3m2d_ca_w_1_120_s_0_140 = 1.37e-04  mcm3m2d_cc_w_1_120_s_0_140 = 1.21e-10  mcm3m2d_cf_w_1_120_s_0_140 = 7.64e-12
+ mcm3m2d_ca_w_1_120_s_0_175 = 1.37e-04  mcm3m2d_cc_w_1_120_s_0_175 = 1.13e-10  mcm3m2d_cf_w_1_120_s_0_175 = 9.75e-12
+ mcm3m2d_ca_w_1_120_s_0_210 = 1.37e-04  mcm3m2d_cc_w_1_120_s_0_210 = 1.06e-10  mcm3m2d_cf_w_1_120_s_0_210 = 1.18e-11
+ mcm3m2d_ca_w_1_120_s_0_280 = 1.37e-04  mcm3m2d_cc_w_1_120_s_0_280 = 8.79e-11  mcm3m2d_cf_w_1_120_s_0_280 = 1.57e-11
+ mcm3m2d_ca_w_1_120_s_0_350 = 1.37e-04  mcm3m2d_cc_w_1_120_s_0_350 = 7.25e-11  mcm3m2d_cf_w_1_120_s_0_350 = 1.94e-11
+ mcm3m2d_ca_w_1_120_s_0_420 = 1.37e-04  mcm3m2d_cc_w_1_120_s_0_420 = 6.00e-11  mcm3m2d_cf_w_1_120_s_0_420 = 2.30e-11
+ mcm3m2d_ca_w_1_120_s_0_560 = 1.37e-04  mcm3m2d_cc_w_1_120_s_0_560 = 4.27e-11  mcm3m2d_cf_w_1_120_s_0_560 = 2.92e-11
+ mcm3m2d_ca_w_1_120_s_0_840 = 1.37e-04  mcm3m2d_cc_w_1_120_s_0_840 = 2.44e-11  mcm3m2d_cf_w_1_120_s_0_840 = 3.88e-11
+ mcm3m2d_ca_w_1_120_s_1_540 = 1.37e-04  mcm3m2d_cc_w_1_120_s_1_540 = 7.57e-12  mcm3m2d_cf_w_1_120_s_1_540 = 5.17e-11
+ mcm3m2d_ca_w_1_120_s_3_500 = 1.37e-04  mcm3m2d_cc_w_1_120_s_3_500 = 4.60e-13  mcm3m2d_cf_w_1_120_s_3_500 = 5.87e-11
+ mcm3m2p1_ca_w_0_140_s_0_140 = 1.44e-04  mcm3m2p1_cc_w_0_140_s_0_140 = 1.09e-10  mcm3m2p1_cf_w_0_140_s_0_140 = 7.98e-12
+ mcm3m2p1_ca_w_0_140_s_0_175 = 1.44e-04  mcm3m2p1_cc_w_0_140_s_0_175 = 1.04e-10  mcm3m2p1_cf_w_0_140_s_0_175 = 1.02e-11
+ mcm3m2p1_ca_w_0_140_s_0_210 = 1.44e-04  mcm3m2p1_cc_w_0_140_s_0_210 = 9.76e-11  mcm3m2p1_cf_w_0_140_s_0_210 = 1.24e-11
+ mcm3m2p1_ca_w_0_140_s_0_280 = 1.44e-04  mcm3m2p1_cc_w_0_140_s_0_280 = 8.08e-11  mcm3m2p1_cf_w_0_140_s_0_280 = 1.65e-11
+ mcm3m2p1_ca_w_0_140_s_0_350 = 1.44e-04  mcm3m2p1_cc_w_0_140_s_0_350 = 6.62e-11  mcm3m2p1_cf_w_0_140_s_0_350 = 2.03e-11
+ mcm3m2p1_ca_w_0_140_s_0_420 = 1.44e-04  mcm3m2p1_cc_w_0_140_s_0_420 = 5.44e-11  mcm3m2p1_cf_w_0_140_s_0_420 = 2.42e-11
+ mcm3m2p1_ca_w_0_140_s_0_560 = 1.44e-04  mcm3m2p1_cc_w_0_140_s_0_560 = 3.80e-11  mcm3m2p1_cf_w_0_140_s_0_560 = 3.05e-11
+ mcm3m2p1_ca_w_0_140_s_0_840 = 1.44e-04  mcm3m2p1_cc_w_0_140_s_0_840 = 2.07e-11  mcm3m2p1_cf_w_0_140_s_0_840 = 4.05e-11
+ mcm3m2p1_ca_w_0_140_s_1_540 = 1.44e-04  mcm3m2p1_cc_w_0_140_s_1_540 = 5.51e-12  mcm3m2p1_cf_w_0_140_s_1_540 = 5.28e-11
+ mcm3m2p1_ca_w_0_140_s_3_500 = 1.44e-04  mcm3m2p1_cc_w_0_140_s_3_500 = 2.00e-13  mcm3m2p1_cf_w_0_140_s_3_500 = 5.81e-11
+ mcm3m2p1_ca_w_1_120_s_0_140 = 1.44e-04  mcm3m2p1_cc_w_1_120_s_0_140 = 1.18e-10  mcm3m2p1_cf_w_1_120_s_0_140 = 8.03e-12
+ mcm3m2p1_ca_w_1_120_s_0_175 = 1.44e-04  mcm3m2p1_cc_w_1_120_s_0_175 = 1.11e-10  mcm3m2p1_cf_w_1_120_s_0_175 = 1.03e-11
+ mcm3m2p1_ca_w_1_120_s_0_210 = 1.44e-04  mcm3m2p1_cc_w_1_120_s_0_210 = 1.03e-10  mcm3m2p1_cf_w_1_120_s_0_210 = 1.24e-11
+ mcm3m2p1_ca_w_1_120_s_0_280 = 1.44e-04  mcm3m2p1_cc_w_1_120_s_0_280 = 8.56e-11  mcm3m2p1_cf_w_1_120_s_0_280 = 1.65e-11
+ mcm3m2p1_ca_w_1_120_s_0_350 = 1.44e-04  mcm3m2p1_cc_w_1_120_s_0_350 = 7.03e-11  mcm3m2p1_cf_w_1_120_s_0_350 = 2.05e-11
+ mcm3m2p1_ca_w_1_120_s_0_420 = 1.44e-04  mcm3m2p1_cc_w_1_120_s_0_420 = 5.76e-11  mcm3m2p1_cf_w_1_120_s_0_420 = 2.42e-11
+ mcm3m2p1_ca_w_1_120_s_0_560 = 1.44e-04  mcm3m2p1_cc_w_1_120_s_0_560 = 4.03e-11  mcm3m2p1_cf_w_1_120_s_0_560 = 3.07e-11
+ mcm3m2p1_ca_w_1_120_s_0_840 = 1.44e-04  mcm3m2p1_cc_w_1_120_s_0_840 = 2.21e-11  mcm3m2p1_cf_w_1_120_s_0_840 = 4.08e-11
+ mcm3m2p1_ca_w_1_120_s_1_540 = 1.44e-04  mcm3m2p1_cc_w_1_120_s_1_540 = 6.04e-12  mcm3m2p1_cf_w_1_120_s_1_540 = 5.35e-11
+ mcm3m2p1_ca_w_1_120_s_3_500 = 1.44e-04  mcm3m2p1_cc_w_1_120_s_3_500 = 2.55e-13  mcm3m2p1_cf_w_1_120_s_3_500 = 5.94e-11
+ mcm3m2l1_ca_w_0_140_s_0_140 = 1.58e-04  mcm3m2l1_cc_w_0_140_s_0_140 = 1.08e-10  mcm3m2l1_cf_w_0_140_s_0_140 = 8.81e-12
+ mcm3m2l1_ca_w_0_140_s_0_175 = 1.58e-04  mcm3m2l1_cc_w_0_140_s_0_175 = 1.03e-10  mcm3m2l1_cf_w_0_140_s_0_175 = 1.13e-11
+ mcm3m2l1_ca_w_0_140_s_0_210 = 1.58e-04  mcm3m2l1_cc_w_0_140_s_0_210 = 9.56e-11  mcm3m2l1_cf_w_0_140_s_0_210 = 1.37e-11
+ mcm3m2l1_ca_w_0_140_s_0_280 = 1.58e-04  mcm3m2l1_cc_w_0_140_s_0_280 = 7.90e-11  mcm3m2l1_cf_w_0_140_s_0_280 = 1.83e-11
+ mcm3m2l1_ca_w_0_140_s_0_350 = 1.58e-04  mcm3m2l1_cc_w_0_140_s_0_350 = 6.40e-11  mcm3m2l1_cf_w_0_140_s_0_350 = 2.27e-11
+ mcm3m2l1_ca_w_0_140_s_0_420 = 1.58e-04  mcm3m2l1_cc_w_0_140_s_0_420 = 5.17e-11  mcm3m2l1_cf_w_0_140_s_0_420 = 2.68e-11
+ mcm3m2l1_ca_w_0_140_s_0_560 = 1.58e-04  mcm3m2l1_cc_w_0_140_s_0_560 = 3.50e-11  mcm3m2l1_cf_w_0_140_s_0_560 = 3.39e-11
+ mcm3m2l1_ca_w_0_140_s_0_840 = 1.58e-04  mcm3m2l1_cc_w_0_140_s_0_840 = 1.77e-11  mcm3m2l1_cf_w_0_140_s_0_840 = 4.46e-11
+ mcm3m2l1_ca_w_0_140_s_1_540 = 1.58e-04  mcm3m2l1_cc_w_0_140_s_1_540 = 3.75e-12  mcm3m2l1_cf_w_0_140_s_1_540 = 5.67e-11
+ mcm3m2l1_ca_w_0_140_s_3_500 = 1.58e-04  mcm3m2l1_cc_w_0_140_s_3_500 = 8.50e-14  mcm3m2l1_cf_w_0_140_s_3_500 = 6.05e-11
+ mcm3m2l1_ca_w_1_120_s_0_140 = 1.58e-04  mcm3m2l1_cc_w_1_120_s_0_140 = 1.13e-10  mcm3m2l1_cf_w_1_120_s_0_140 = 8.84e-12
+ mcm3m2l1_ca_w_1_120_s_0_175 = 1.58e-04  mcm3m2l1_cc_w_1_120_s_0_175 = 1.07e-10  mcm3m2l1_cf_w_1_120_s_0_175 = 1.13e-11
+ mcm3m2l1_ca_w_1_120_s_0_210 = 1.58e-04  mcm3m2l1_cc_w_1_120_s_0_210 = 9.90e-11  mcm3m2l1_cf_w_1_120_s_0_210 = 1.37e-11
+ mcm3m2l1_ca_w_1_120_s_0_280 = 1.58e-04  mcm3m2l1_cc_w_1_120_s_0_280 = 8.15e-11  mcm3m2l1_cf_w_1_120_s_0_280 = 1.83e-11
+ mcm3m2l1_ca_w_1_120_s_0_350 = 1.58e-04  mcm3m2l1_cc_w_1_120_s_0_350 = 6.62e-11  mcm3m2l1_cf_w_1_120_s_0_350 = 2.27e-11
+ mcm3m2l1_ca_w_1_120_s_0_420 = 1.58e-04  mcm3m2l1_cc_w_1_120_s_0_420 = 5.37e-11  mcm3m2l1_cf_w_1_120_s_0_420 = 2.68e-11
+ mcm3m2l1_ca_w_1_120_s_0_560 = 1.58e-04  mcm3m2l1_cc_w_1_120_s_0_560 = 3.63e-11  mcm3m2l1_cf_w_1_120_s_0_560 = 3.41e-11
+ mcm3m2l1_ca_w_1_120_s_0_840 = 1.58e-04  mcm3m2l1_cc_w_1_120_s_0_840 = 1.84e-11  mcm3m2l1_cf_w_1_120_s_0_840 = 4.49e-11
+ mcm3m2l1_ca_w_1_120_s_1_540 = 1.58e-04  mcm3m2l1_cc_w_1_120_s_1_540 = 3.93e-12  mcm3m2l1_cf_w_1_120_s_1_540 = 5.71e-11
+ mcm3m2l1_ca_w_1_120_s_3_500 = 1.58e-04  mcm3m2l1_cc_w_1_120_s_3_500 = 1.10e-13  mcm3m2l1_cf_w_1_120_s_3_500 = 6.13e-11
+ mcm3m2m1_ca_w_0_140_s_0_140 = 3.31e-04  mcm3m2m1_cc_w_0_140_s_0_140 = 9.50e-11  mcm3m2m1_cf_w_0_140_s_0_140 = 1.76e-11
+ mcm3m2m1_ca_w_0_140_s_0_175 = 3.31e-04  mcm3m2m1_cc_w_0_140_s_0_175 = 8.95e-11  mcm3m2m1_cf_w_0_140_s_0_175 = 2.30e-11
+ mcm3m2m1_ca_w_0_140_s_0_210 = 3.31e-04  mcm3m2m1_cc_w_0_140_s_0_210 = 8.16e-11  mcm3m2m1_cf_w_0_140_s_0_210 = 2.82e-11
+ mcm3m2m1_ca_w_0_140_s_0_280 = 3.31e-04  mcm3m2m1_cc_w_0_140_s_0_280 = 6.45e-11  mcm3m2m1_cf_w_0_140_s_0_280 = 3.75e-11
+ mcm3m2m1_ca_w_0_140_s_0_350 = 3.31e-04  mcm3m2m1_cc_w_0_140_s_0_350 = 4.92e-11  mcm3m2m1_cf_w_0_140_s_0_350 = 4.58e-11
+ mcm3m2m1_ca_w_0_140_s_0_420 = 3.31e-04  mcm3m2m1_cc_w_0_140_s_0_420 = 3.72e-11  mcm3m2m1_cf_w_0_140_s_0_420 = 5.31e-11
+ mcm3m2m1_ca_w_0_140_s_0_560 = 3.31e-04  mcm3m2m1_cc_w_0_140_s_0_560 = 2.16e-11  mcm3m2m1_cf_w_0_140_s_0_560 = 6.43e-11
+ mcm3m2m1_ca_w_0_140_s_0_840 = 3.31e-04  mcm3m2m1_cc_w_0_140_s_0_840 = 7.62e-12  mcm3m2m1_cf_w_0_140_s_0_840 = 7.71e-11
+ mcm3m2m1_ca_w_0_140_s_1_540 = 3.31e-04  mcm3m2m1_cc_w_0_140_s_1_540 = 7.25e-13  mcm3m2m1_cf_w_0_140_s_1_540 = 8.52e-11
+ mcm3m2m1_ca_w_0_140_s_3_500 = 3.31e-04  mcm3m2m1_cc_w_0_140_s_3_500 = 2.50e-14  mcm3m2m1_cf_w_0_140_s_3_500 = 8.69e-11
+ mcm3m2m1_ca_w_1_120_s_0_140 = 3.31e-04  mcm3m2m1_cc_w_1_120_s_0_140 = 9.70e-11  mcm3m2m1_cf_w_1_120_s_0_140 = 1.76e-11
+ mcm3m2m1_ca_w_1_120_s_0_175 = 3.31e-04  mcm3m2m1_cc_w_1_120_s_0_175 = 9.06e-11  mcm3m2m1_cf_w_1_120_s_0_175 = 2.30e-11
+ mcm3m2m1_ca_w_1_120_s_0_210 = 3.31e-04  mcm3m2m1_cc_w_1_120_s_0_210 = 8.26e-11  mcm3m2m1_cf_w_1_120_s_0_210 = 2.81e-11
+ mcm3m2m1_ca_w_1_120_s_0_280 = 3.31e-04  mcm3m2m1_cc_w_1_120_s_0_280 = 6.50e-11  mcm3m2m1_cf_w_1_120_s_0_280 = 3.75e-11
+ mcm3m2m1_ca_w_1_120_s_0_350 = 3.31e-04  mcm3m2m1_cc_w_1_120_s_0_350 = 4.98e-11  mcm3m2m1_cf_w_1_120_s_0_350 = 4.58e-11
+ mcm3m2m1_ca_w_1_120_s_0_420 = 3.31e-04  mcm3m2m1_cc_w_1_120_s_0_420 = 3.76e-11  mcm3m2m1_cf_w_1_120_s_0_420 = 5.32e-11
+ mcm3m2m1_ca_w_1_120_s_0_560 = 3.31e-04  mcm3m2m1_cc_w_1_120_s_0_560 = 2.20e-11  mcm3m2m1_cf_w_1_120_s_0_560 = 6.45e-11
+ mcm3m2m1_ca_w_1_120_s_0_840 = 3.31e-04  mcm3m2m1_cc_w_1_120_s_0_840 = 7.70e-12  mcm3m2m1_cf_w_1_120_s_0_840 = 7.72e-11
+ mcm3m2m1_ca_w_1_120_s_1_540 = 3.31e-04  mcm3m2m1_cc_w_1_120_s_1_540 = 7.00e-13  mcm3m2m1_cf_w_1_120_s_1_540 = 8.54e-11
+ mcm3m2m1_ca_w_1_120_s_3_500 = 3.31e-04  mcm3m2m1_cc_w_1_120_s_3_500 = 5.00e-14  mcm3m2m1_cf_w_1_120_s_3_500 = 8.70e-11
+ mcm4m2f_ca_w_0_140_s_0_140 = 4.50e-05  mcm4m2f_cc_w_0_140_s_0_140 = 1.20e-10  mcm4m2f_cf_w_0_140_s_0_140 = 2.64e-12
+ mcm4m2f_ca_w_0_140_s_0_175 = 4.50e-05  mcm4m2f_cc_w_0_140_s_0_175 = 1.15e-10  mcm4m2f_cf_w_0_140_s_0_175 = 3.41e-12
+ mcm4m2f_ca_w_0_140_s_0_210 = 4.50e-05  mcm4m2f_cc_w_0_140_s_0_210 = 1.09e-10  mcm4m2f_cf_w_0_140_s_0_210 = 4.20e-12
+ mcm4m2f_ca_w_0_140_s_0_280 = 4.50e-05  mcm4m2f_cc_w_0_140_s_0_280 = 9.33e-11  mcm4m2f_cf_w_0_140_s_0_280 = 5.71e-12
+ mcm4m2f_ca_w_0_140_s_0_350 = 4.50e-05  mcm4m2f_cc_w_0_140_s_0_350 = 8.01e-11  mcm4m2f_cf_w_0_140_s_0_350 = 7.20e-12
+ mcm4m2f_ca_w_0_140_s_0_420 = 4.50e-05  mcm4m2f_cc_w_0_140_s_0_420 = 6.82e-11  mcm4m2f_cf_w_0_140_s_0_420 = 8.73e-12
+ mcm4m2f_ca_w_0_140_s_0_560 = 4.50e-05  mcm4m2f_cc_w_0_140_s_0_560 = 5.27e-11  mcm4m2f_cf_w_0_140_s_0_560 = 1.15e-11
+ mcm4m2f_ca_w_0_140_s_0_840 = 4.50e-05  mcm4m2f_cc_w_0_140_s_0_840 = 3.54e-11  mcm4m2f_cf_w_0_140_s_0_840 = 1.67e-11
+ mcm4m2f_ca_w_0_140_s_1_540 = 4.50e-05  mcm4m2f_cc_w_0_140_s_1_540 = 1.65e-11  mcm4m2f_cf_w_0_140_s_1_540 = 2.66e-11
+ mcm4m2f_ca_w_0_140_s_3_500 = 4.50e-05  mcm4m2f_cc_w_0_140_s_3_500 = 2.70e-12  mcm4m2f_cf_w_0_140_s_3_500 = 3.77e-11
+ mcm4m2f_ca_w_1_120_s_0_140 = 4.50e-05  mcm4m2f_cc_w_1_120_s_0_140 = 1.37e-10  mcm4m2f_cf_w_1_120_s_0_140 = 2.67e-12
+ mcm4m2f_ca_w_1_120_s_0_175 = 4.50e-05  mcm4m2f_cc_w_1_120_s_0_175 = 1.31e-10  mcm4m2f_cf_w_1_120_s_0_175 = 3.45e-12
+ mcm4m2f_ca_w_1_120_s_0_210 = 4.50e-05  mcm4m2f_cc_w_1_120_s_0_210 = 1.24e-10  mcm4m2f_cf_w_1_120_s_0_210 = 4.23e-12
+ mcm4m2f_ca_w_1_120_s_0_280 = 4.50e-05  mcm4m2f_cc_w_1_120_s_0_280 = 1.06e-10  mcm4m2f_cf_w_1_120_s_0_280 = 5.74e-12
+ mcm4m2f_ca_w_1_120_s_0_350 = 4.50e-05  mcm4m2f_cc_w_1_120_s_0_350 = 9.04e-11  mcm4m2f_cf_w_1_120_s_0_350 = 7.25e-12
+ mcm4m2f_ca_w_1_120_s_0_420 = 4.50e-05  mcm4m2f_cc_w_1_120_s_0_420 = 7.77e-11  mcm4m2f_cf_w_1_120_s_0_420 = 8.73e-12
+ mcm4m2f_ca_w_1_120_s_0_560 = 4.50e-05  mcm4m2f_cc_w_1_120_s_0_560 = 6.01e-11  mcm4m2f_cf_w_1_120_s_0_560 = 1.16e-11
+ mcm4m2f_ca_w_1_120_s_0_840 = 4.50e-05  mcm4m2f_cc_w_1_120_s_0_840 = 4.05e-11  mcm4m2f_cf_w_1_120_s_0_840 = 1.69e-11
+ mcm4m2f_ca_w_1_120_s_1_540 = 4.50e-05  mcm4m2f_cc_w_1_120_s_1_540 = 1.90e-11  mcm4m2f_cf_w_1_120_s_1_540 = 2.72e-11
+ mcm4m2f_ca_w_1_120_s_3_500 = 4.50e-05  mcm4m2f_cc_w_1_120_s_3_500 = 3.18e-12  mcm4m2f_cf_w_1_120_s_3_500 = 3.97e-11
+ mcm4m2d_ca_w_0_140_s_0_140 = 4.87e-05  mcm4m2d_cc_w_0_140_s_0_140 = 1.20e-10  mcm4m2d_cf_w_0_140_s_0_140 = 2.86e-12
+ mcm4m2d_ca_w_0_140_s_0_175 = 4.87e-05  mcm4m2d_cc_w_0_140_s_0_175 = 1.15e-10  mcm4m2d_cf_w_0_140_s_0_175 = 3.69e-12
+ mcm4m2d_ca_w_0_140_s_0_210 = 4.87e-05  mcm4m2d_cc_w_0_140_s_0_210 = 1.08e-10  mcm4m2d_cf_w_0_140_s_0_210 = 4.54e-12
+ mcm4m2d_ca_w_0_140_s_0_280 = 4.87e-05  mcm4m2d_cc_w_0_140_s_0_280 = 9.27e-11  mcm4m2d_cf_w_0_140_s_0_280 = 6.18e-12
+ mcm4m2d_ca_w_0_140_s_0_350 = 4.87e-05  mcm4m2d_cc_w_0_140_s_0_350 = 7.94e-11  mcm4m2d_cf_w_0_140_s_0_350 = 7.79e-12
+ mcm4m2d_ca_w_0_140_s_0_420 = 4.87e-05  mcm4m2d_cc_w_0_140_s_0_420 = 6.74e-11  mcm4m2d_cf_w_0_140_s_0_420 = 9.42e-12
+ mcm4m2d_ca_w_0_140_s_0_560 = 4.87e-05  mcm4m2d_cc_w_0_140_s_0_560 = 5.16e-11  mcm4m2d_cf_w_0_140_s_0_560 = 1.24e-11
+ mcm4m2d_ca_w_0_140_s_0_840 = 4.87e-05  mcm4m2d_cc_w_0_140_s_0_840 = 3.44e-11  mcm4m2d_cf_w_0_140_s_0_840 = 1.79e-11
+ mcm4m2d_ca_w_0_140_s_1_540 = 4.87e-05  mcm4m2d_cc_w_0_140_s_1_540 = 1.54e-11  mcm4m2d_cf_w_0_140_s_1_540 = 2.82e-11
+ mcm4m2d_ca_w_0_140_s_3_500 = 4.87e-05  mcm4m2d_cc_w_0_140_s_3_500 = 2.21e-12  mcm4m2d_cf_w_0_140_s_3_500 = 3.92e-11
+ mcm4m2d_ca_w_1_120_s_0_140 = 4.87e-05  mcm4m2d_cc_w_1_120_s_0_140 = 1.36e-10  mcm4m2d_cf_w_1_120_s_0_140 = 2.90e-12
+ mcm4m2d_ca_w_1_120_s_0_175 = 4.87e-05  mcm4m2d_cc_w_1_120_s_0_175 = 1.30e-10  mcm4m2d_cf_w_1_120_s_0_175 = 3.73e-12
+ mcm4m2d_ca_w_1_120_s_0_210 = 4.87e-05  mcm4m2d_cc_w_1_120_s_0_210 = 1.22e-10  mcm4m2d_cf_w_1_120_s_0_210 = 4.56e-12
+ mcm4m2d_ca_w_1_120_s_0_280 = 4.87e-05  mcm4m2d_cc_w_1_120_s_0_280 = 1.05e-10  mcm4m2d_cf_w_1_120_s_0_280 = 6.21e-12
+ mcm4m2d_ca_w_1_120_s_0_350 = 4.87e-05  mcm4m2d_cc_w_1_120_s_0_350 = 8.88e-11  mcm4m2d_cf_w_1_120_s_0_350 = 7.83e-12
+ mcm4m2d_ca_w_1_120_s_0_420 = 4.87e-05  mcm4m2d_cc_w_1_120_s_0_420 = 7.61e-11  mcm4m2d_cf_w_1_120_s_0_420 = 9.43e-12
+ mcm4m2d_ca_w_1_120_s_0_560 = 4.87e-05  mcm4m2d_cc_w_1_120_s_0_560 = 5.84e-11  mcm4m2d_cf_w_1_120_s_0_560 = 1.25e-11
+ mcm4m2d_ca_w_1_120_s_0_840 = 4.87e-05  mcm4m2d_cc_w_1_120_s_0_840 = 3.88e-11  mcm4m2d_cf_w_1_120_s_0_840 = 1.82e-11
+ mcm4m2d_ca_w_1_120_s_1_540 = 4.87e-05  mcm4m2d_cc_w_1_120_s_1_540 = 1.76e-11  mcm4m2d_cf_w_1_120_s_1_540 = 2.90e-11
+ mcm4m2d_ca_w_1_120_s_3_500 = 4.87e-05  mcm4m2d_cc_w_1_120_s_3_500 = 2.57e-12  mcm4m2d_cf_w_1_120_s_3_500 = 4.11e-11
+ mcm4m2p1_ca_w_0_140_s_0_140 = 5.50e-05  mcm4m2p1_cc_w_0_140_s_0_140 = 1.18e-10  mcm4m2p1_cf_w_0_140_s_0_140 = 3.23e-12
+ mcm4m2p1_ca_w_0_140_s_0_175 = 5.50e-05  mcm4m2p1_cc_w_0_140_s_0_175 = 1.14e-10  mcm4m2p1_cf_w_0_140_s_0_175 = 4.17e-12
+ mcm4m2p1_ca_w_0_140_s_0_210 = 5.50e-05  mcm4m2p1_cc_w_0_140_s_0_210 = 1.08e-10  mcm4m2p1_cf_w_0_140_s_0_210 = 5.14e-12
+ mcm4m2p1_ca_w_0_140_s_0_280 = 5.50e-05  mcm4m2p1_cc_w_0_140_s_0_280 = 9.16e-11  mcm4m2p1_cf_w_0_140_s_0_280 = 6.99e-12
+ mcm4m2p1_ca_w_0_140_s_0_350 = 5.50e-05  mcm4m2p1_cc_w_0_140_s_0_350 = 7.76e-11  mcm4m2p1_cf_w_0_140_s_0_350 = 8.78e-12
+ mcm4m2p1_ca_w_0_140_s_0_420 = 5.50e-05  mcm4m2p1_cc_w_0_140_s_0_420 = 6.59e-11  mcm4m2p1_cf_w_0_140_s_0_420 = 1.06e-11
+ mcm4m2p1_ca_w_0_140_s_0_560 = 5.50e-05  mcm4m2p1_cc_w_0_140_s_0_560 = 5.03e-11  mcm4m2p1_cf_w_0_140_s_0_560 = 1.40e-11
+ mcm4m2p1_ca_w_0_140_s_0_840 = 5.50e-05  mcm4m2p1_cc_w_0_140_s_0_840 = 3.26e-11  mcm4m2p1_cf_w_0_140_s_0_840 = 2.00e-11
+ mcm4m2p1_ca_w_0_140_s_1_540 = 5.50e-05  mcm4m2p1_cc_w_0_140_s_1_540 = 1.38e-11  mcm4m2p1_cf_w_0_140_s_1_540 = 3.10e-11
+ mcm4m2p1_ca_w_0_140_s_3_500 = 5.50e-05  mcm4m2p1_cc_w_0_140_s_3_500 = 1.65e-12  mcm4m2p1_cf_w_0_140_s_3_500 = 4.14e-11
+ mcm4m2p1_ca_w_1_120_s_0_140 = 5.50e-05  mcm4m2p1_cc_w_1_120_s_0_140 = 1.34e-10  mcm4m2p1_cf_w_1_120_s_0_140 = 3.31e-12
+ mcm4m2p1_ca_w_1_120_s_0_175 = 5.50e-05  mcm4m2p1_cc_w_1_120_s_0_175 = 1.27e-10  mcm4m2p1_cf_w_1_120_s_0_175 = 4.26e-12
+ mcm4m2p1_ca_w_1_120_s_0_210 = 5.50e-05  mcm4m2p1_cc_w_1_120_s_0_210 = 1.20e-10  mcm4m2p1_cf_w_1_120_s_0_210 = 5.20e-12
+ mcm4m2p1_ca_w_1_120_s_0_280 = 5.50e-05  mcm4m2p1_cc_w_1_120_s_0_280 = 1.02e-10  mcm4m2p1_cf_w_1_120_s_0_280 = 7.04e-12
+ mcm4m2p1_ca_w_1_120_s_0_350 = 5.50e-05  mcm4m2p1_cc_w_1_120_s_0_350 = 8.63e-11  mcm4m2p1_cf_w_1_120_s_0_350 = 8.86e-12
+ mcm4m2p1_ca_w_1_120_s_0_420 = 5.50e-05  mcm4m2p1_cc_w_1_120_s_0_420 = 7.36e-11  mcm4m2p1_cf_w_1_120_s_0_420 = 1.07e-11
+ mcm4m2p1_ca_w_1_120_s_0_560 = 5.50e-05  mcm4m2p1_cc_w_1_120_s_0_560 = 5.59e-11  mcm4m2p1_cf_w_1_120_s_0_560 = 1.41e-11
+ mcm4m2p1_ca_w_1_120_s_0_840 = 5.50e-05  mcm4m2p1_cc_w_1_120_s_0_840 = 3.63e-11  mcm4m2p1_cf_w_1_120_s_0_840 = 2.03e-11
+ mcm4m2p1_ca_w_1_120_s_1_540 = 5.50e-05  mcm4m2p1_cc_w_1_120_s_1_540 = 1.55e-11  mcm4m2p1_cf_w_1_120_s_1_540 = 3.18e-11
+ mcm4m2p1_ca_w_1_120_s_3_500 = 5.50e-05  mcm4m2p1_cc_w_1_120_s_3_500 = 1.90e-12  mcm4m2p1_cf_w_1_120_s_3_500 = 4.33e-11
+ mcm4m2l1_ca_w_0_140_s_0_140 = 6.98e-05  mcm4m2l1_cc_w_0_140_s_0_140 = 1.16e-10  mcm4m2l1_cf_w_0_140_s_0_140 = 4.06e-12
+ mcm4m2l1_ca_w_0_140_s_0_175 = 6.98e-05  mcm4m2l1_cc_w_0_140_s_0_175 = 1.12e-10  mcm4m2l1_cf_w_0_140_s_0_175 = 5.25e-12
+ mcm4m2l1_ca_w_0_140_s_0_210 = 6.98e-05  mcm4m2l1_cc_w_0_140_s_0_210 = 1.05e-10  mcm4m2l1_cf_w_0_140_s_0_210 = 6.46e-12
+ mcm4m2l1_ca_w_0_140_s_0_280 = 6.98e-05  mcm4m2l1_cc_w_0_140_s_0_280 = 9.01e-11  mcm4m2l1_cf_w_0_140_s_0_280 = 8.79e-12
+ mcm4m2l1_ca_w_0_140_s_0_350 = 6.98e-05  mcm4m2l1_cc_w_0_140_s_0_350 = 7.55e-11  mcm4m2l1_cf_w_0_140_s_0_350 = 1.11e-11
+ mcm4m2l1_ca_w_0_140_s_0_420 = 6.98e-05  mcm4m2l1_cc_w_0_140_s_0_420 = 6.36e-11  mcm4m2l1_cf_w_0_140_s_0_420 = 1.33e-11
+ mcm4m2l1_ca_w_0_140_s_0_560 = 6.98e-05  mcm4m2l1_cc_w_0_140_s_0_560 = 4.73e-11  mcm4m2l1_cf_w_0_140_s_0_560 = 1.75e-11
+ mcm4m2l1_ca_w_0_140_s_0_840 = 6.98e-05  mcm4m2l1_cc_w_0_140_s_0_840 = 2.93e-11  mcm4m2l1_cf_w_0_140_s_0_840 = 2.47e-11
+ mcm4m2l1_ca_w_0_140_s_1_540 = 6.98e-05  mcm4m2l1_cc_w_0_140_s_1_540 = 1.11e-11  mcm4m2l1_cf_w_0_140_s_1_540 = 3.66e-11
+ mcm4m2l1_ca_w_0_140_s_3_500 = 6.98e-05  mcm4m2l1_cc_w_0_140_s_3_500 = 1.01e-12  mcm4m2l1_cf_w_0_140_s_3_500 = 4.56e-11
+ mcm4m2l1_ca_w_1_120_s_0_140 = 6.98e-05  mcm4m2l1_cc_w_1_120_s_0_140 = 1.31e-10  mcm4m2l1_cf_w_1_120_s_0_140 = 4.10e-12
+ mcm4m2l1_ca_w_1_120_s_0_175 = 6.98e-05  mcm4m2l1_cc_w_1_120_s_0_175 = 1.24e-10  mcm4m2l1_cf_w_1_120_s_0_175 = 5.30e-12
+ mcm4m2l1_ca_w_1_120_s_0_210 = 6.98e-05  mcm4m2l1_cc_w_1_120_s_0_210 = 1.16e-10  mcm4m2l1_cf_w_1_120_s_0_210 = 6.49e-12
+ mcm4m2l1_ca_w_1_120_s_0_280 = 6.98e-05  mcm4m2l1_cc_w_1_120_s_0_280 = 9.77e-11  mcm4m2l1_cf_w_1_120_s_0_280 = 8.83e-12
+ mcm4m2l1_ca_w_1_120_s_0_350 = 6.98e-05  mcm4m2l1_cc_w_1_120_s_0_350 = 8.23e-11  mcm4m2l1_cf_w_1_120_s_0_350 = 1.11e-11
+ mcm4m2l1_ca_w_1_120_s_0_420 = 6.98e-05  mcm4m2l1_cc_w_1_120_s_0_420 = 6.98e-11  mcm4m2l1_cf_w_1_120_s_0_420 = 1.33e-11
+ mcm4m2l1_ca_w_1_120_s_0_560 = 6.98e-05  mcm4m2l1_cc_w_1_120_s_0_560 = 5.18e-11  mcm4m2l1_cf_w_1_120_s_0_560 = 1.75e-11
+ mcm4m2l1_ca_w_1_120_s_0_840 = 6.98e-05  mcm4m2l1_cc_w_1_120_s_0_840 = 3.24e-11  mcm4m2l1_cf_w_1_120_s_0_840 = 2.50e-11
+ mcm4m2l1_ca_w_1_120_s_1_540 = 6.98e-05  mcm4m2l1_cc_w_1_120_s_1_540 = 1.24e-11  mcm4m2l1_cf_w_1_120_s_1_540 = 3.74e-11
+ mcm4m2l1_ca_w_1_120_s_3_500 = 6.98e-05  mcm4m2l1_cc_w_1_120_s_3_500 = 1.14e-12  mcm4m2l1_cf_w_1_120_s_3_500 = 4.76e-11
+ mcm4m2m1_ca_w_0_140_s_0_140 = 2.42e-04  mcm4m2m1_cc_w_0_140_s_0_140 = 1.05e-10  mcm4m2m1_cf_w_0_140_s_0_140 = 1.28e-11
+ mcm4m2m1_ca_w_0_140_s_0_175 = 2.42e-04  mcm4m2m1_cc_w_0_140_s_0_175 = 9.87e-11  mcm4m2m1_cf_w_0_140_s_0_175 = 1.70e-11
+ mcm4m2m1_ca_w_0_140_s_0_210 = 2.42e-04  mcm4m2m1_cc_w_0_140_s_0_210 = 9.11e-11  mcm4m2m1_cf_w_0_140_s_0_210 = 2.09e-11
+ mcm4m2m1_ca_w_0_140_s_0_280 = 2.42e-04  mcm4m2m1_cc_w_0_140_s_0_280 = 7.51e-11  mcm4m2m1_cf_w_0_140_s_0_280 = 2.80e-11
+ mcm4m2m1_ca_w_0_140_s_0_350 = 2.42e-04  mcm4m2m1_cc_w_0_140_s_0_350 = 6.06e-11  mcm4m2m1_cf_w_0_140_s_0_350 = 3.43e-11
+ mcm4m2m1_ca_w_0_140_s_0_420 = 2.42e-04  mcm4m2m1_cc_w_0_140_s_0_420 = 4.86e-11  mcm4m2m1_cf_w_0_140_s_0_420 = 3.97e-11
+ mcm4m2m1_ca_w_0_140_s_0_560 = 2.42e-04  mcm4m2m1_cc_w_0_140_s_0_560 = 3.31e-11  mcm4m2m1_cf_w_0_140_s_0_560 = 4.86e-11
+ mcm4m2m1_ca_w_0_140_s_0_840 = 2.42e-04  mcm4m2m1_cc_w_0_140_s_0_840 = 1.74e-11  mcm4m2m1_cf_w_0_140_s_0_840 = 6.05e-11
+ mcm4m2m1_ca_w_0_140_s_1_540 = 2.42e-04  mcm4m2m1_cc_w_0_140_s_1_540 = 4.53e-12  mcm4m2m1_cf_w_0_140_s_1_540 = 7.25e-11
+ mcm4m2m1_ca_w_0_140_s_3_500 = 2.42e-04  mcm4m2m1_cc_w_0_140_s_3_500 = 2.50e-13  mcm4m2m1_cf_w_0_140_s_3_500 = 7.76e-11
+ mcm4m2m1_ca_w_1_120_s_0_140 = 2.42e-04  mcm4m2m1_cc_w_1_120_s_0_140 = 1.13e-10  mcm4m2m1_cf_w_1_120_s_0_140 = 1.28e-11
+ mcm4m2m1_ca_w_1_120_s_0_175 = 2.42e-04  mcm4m2m1_cc_w_1_120_s_0_175 = 1.07e-10  mcm4m2m1_cf_w_1_120_s_0_175 = 1.70e-11
+ mcm4m2m1_ca_w_1_120_s_0_210 = 2.42e-04  mcm4m2m1_cc_w_1_120_s_0_210 = 9.86e-11  mcm4m2m1_cf_w_1_120_s_0_210 = 2.09e-11
+ mcm4m2m1_ca_w_1_120_s_0_280 = 2.42e-04  mcm4m2m1_cc_w_1_120_s_0_280 = 8.11e-11  mcm4m2m1_cf_w_1_120_s_0_280 = 2.80e-11
+ mcm4m2m1_ca_w_1_120_s_0_350 = 2.42e-04  mcm4m2m1_cc_w_1_120_s_0_350 = 6.57e-11  mcm4m2m1_cf_w_1_120_s_0_350 = 3.43e-11
+ mcm4m2m1_ca_w_1_120_s_0_420 = 2.42e-04  mcm4m2m1_cc_w_1_120_s_0_420 = 5.36e-11  mcm4m2m1_cf_w_1_120_s_0_420 = 3.97e-11
+ mcm4m2m1_ca_w_1_120_s_0_560 = 2.42e-04  mcm4m2m1_cc_w_1_120_s_0_560 = 3.70e-11  mcm4m2m1_cf_w_1_120_s_0_560 = 4.87e-11
+ mcm4m2m1_ca_w_1_120_s_0_840 = 2.42e-04  mcm4m2m1_cc_w_1_120_s_0_840 = 1.99e-11  mcm4m2m1_cf_w_1_120_s_0_840 = 6.07e-11
+ mcm4m2m1_ca_w_1_120_s_1_540 = 2.42e-04  mcm4m2m1_cc_w_1_120_s_1_540 = 5.55e-12  mcm4m2m1_cf_w_1_120_s_1_540 = 7.39e-11
+ mcm4m2m1_ca_w_1_120_s_3_500 = 2.42e-04  mcm4m2m1_cc_w_1_120_s_3_500 = 3.05e-13  mcm4m2m1_cf_w_1_120_s_3_500 = 7.99e-11
+ mcm5m2f_ca_w_0_140_s_0_140 = 3.40e-05  mcm5m2f_cc_w_0_140_s_0_140 = 1.21e-10  mcm5m2f_cf_w_0_140_s_0_140 = 2.00e-12
+ mcm5m2f_ca_w_0_140_s_0_175 = 3.40e-05  mcm5m2f_cc_w_0_140_s_0_175 = 1.17e-10  mcm5m2f_cf_w_0_140_s_0_175 = 2.59e-12
+ mcm5m2f_ca_w_0_140_s_0_210 = 3.40e-05  mcm5m2f_cc_w_0_140_s_0_210 = 1.10e-10  mcm5m2f_cf_w_0_140_s_0_210 = 3.19e-12
+ mcm5m2f_ca_w_0_140_s_0_280 = 3.40e-05  mcm5m2f_cc_w_0_140_s_0_280 = 9.46e-11  mcm5m2f_cf_w_0_140_s_0_280 = 4.35e-12
+ mcm5m2f_ca_w_0_140_s_0_350 = 3.40e-05  mcm5m2f_cc_w_0_140_s_0_350 = 8.24e-11  mcm5m2f_cf_w_0_140_s_0_350 = 5.50e-12
+ mcm5m2f_ca_w_0_140_s_0_420 = 3.40e-05  mcm5m2f_cc_w_0_140_s_0_420 = 7.07e-11  mcm5m2f_cf_w_0_140_s_0_420 = 6.68e-12
+ mcm5m2f_ca_w_0_140_s_0_560 = 3.40e-05  mcm5m2f_cc_w_0_140_s_0_560 = 5.54e-11  mcm5m2f_cf_w_0_140_s_0_560 = 8.86e-12
+ mcm5m2f_ca_w_0_140_s_0_840 = 3.40e-05  mcm5m2f_cc_w_0_140_s_0_840 = 3.90e-11  mcm5m2f_cf_w_0_140_s_0_840 = 1.29e-11
+ mcm5m2f_ca_w_0_140_s_1_540 = 3.40e-05  mcm5m2f_cc_w_0_140_s_1_540 = 2.04e-11  mcm5m2f_cf_w_0_140_s_1_540 = 2.13e-11
+ mcm5m2f_ca_w_0_140_s_3_500 = 3.40e-05  mcm5m2f_cc_w_0_140_s_3_500 = 4.87e-12  mcm5m2f_cf_w_0_140_s_3_500 = 3.28e-11
+ mcm5m2f_ca_w_1_120_s_0_140 = 3.40e-05  mcm5m2f_cc_w_1_120_s_0_140 = 1.41e-10  mcm5m2f_cf_w_1_120_s_0_140 = 2.04e-12
+ mcm5m2f_ca_w_1_120_s_0_175 = 3.40e-05  mcm5m2f_cc_w_1_120_s_0_175 = 1.36e-10  mcm5m2f_cf_w_1_120_s_0_175 = 2.63e-12
+ mcm5m2f_ca_w_1_120_s_0_210 = 3.40e-05  mcm5m2f_cc_w_1_120_s_0_210 = 1.29e-10  mcm5m2f_cf_w_1_120_s_0_210 = 3.22e-12
+ mcm5m2f_ca_w_1_120_s_0_280 = 3.40e-05  mcm5m2f_cc_w_1_120_s_0_280 = 1.11e-10  mcm5m2f_cf_w_1_120_s_0_280 = 4.39e-12
+ mcm5m2f_ca_w_1_120_s_0_350 = 3.40e-05  mcm5m2f_cc_w_1_120_s_0_350 = 9.56e-11  mcm5m2f_cf_w_1_120_s_0_350 = 5.55e-12
+ mcm5m2f_ca_w_1_120_s_0_420 = 3.40e-05  mcm5m2f_cc_w_1_120_s_0_420 = 8.30e-11  mcm5m2f_cf_w_1_120_s_0_420 = 6.68e-12
+ mcm5m2f_ca_w_1_120_s_0_560 = 3.40e-05  mcm5m2f_cc_w_1_120_s_0_560 = 6.53e-11  mcm5m2f_cf_w_1_120_s_0_560 = 8.90e-12
+ mcm5m2f_ca_w_1_120_s_0_840 = 3.40e-05  mcm5m2f_cc_w_1_120_s_0_840 = 4.60e-11  mcm5m2f_cf_w_1_120_s_0_840 = 1.31e-11
+ mcm5m2f_ca_w_1_120_s_1_540 = 3.40e-05  mcm5m2f_cc_w_1_120_s_1_540 = 2.44e-11  mcm5m2f_cf_w_1_120_s_1_540 = 2.18e-11
+ mcm5m2f_ca_w_1_120_s_3_500 = 3.40e-05  mcm5m2f_cc_w_1_120_s_3_500 = 5.97e-12  mcm5m2f_cf_w_1_120_s_3_500 = 3.48e-11
+ mcm5m2d_ca_w_0_140_s_0_140 = 3.77e-05  mcm5m2d_cc_w_0_140_s_0_140 = 1.21e-10  mcm5m2d_cf_w_0_140_s_0_140 = 2.22e-12
+ mcm5m2d_ca_w_0_140_s_0_175 = 3.77e-05  mcm5m2d_cc_w_0_140_s_0_175 = 1.16e-10  mcm5m2d_cf_w_0_140_s_0_175 = 2.87e-12
+ mcm5m2d_ca_w_0_140_s_0_210 = 3.77e-05  mcm5m2d_cc_w_0_140_s_0_210 = 1.10e-10  mcm5m2d_cf_w_0_140_s_0_210 = 3.53e-12
+ mcm5m2d_ca_w_0_140_s_0_280 = 3.77e-05  mcm5m2d_cc_w_0_140_s_0_280 = 9.48e-11  mcm5m2d_cf_w_0_140_s_0_280 = 4.82e-12
+ mcm5m2d_ca_w_0_140_s_0_350 = 3.77e-05  mcm5m2d_cc_w_0_140_s_0_350 = 8.13e-11  mcm5m2d_cf_w_0_140_s_0_350 = 6.07e-12
+ mcm5m2d_ca_w_0_140_s_0_420 = 3.77e-05  mcm5m2d_cc_w_0_140_s_0_420 = 7.00e-11  mcm5m2d_cf_w_0_140_s_0_420 = 7.39e-12
+ mcm5m2d_ca_w_0_140_s_0_560 = 3.77e-05  mcm5m2d_cc_w_0_140_s_0_560 = 5.44e-11  mcm5m2d_cf_w_0_140_s_0_560 = 9.78e-12
+ mcm5m2d_ca_w_0_140_s_0_840 = 3.77e-05  mcm5m2d_cc_w_0_140_s_0_840 = 3.78e-11  mcm5m2d_cf_w_0_140_s_0_840 = 1.42e-11
+ mcm5m2d_ca_w_0_140_s_1_540 = 3.77e-05  mcm5m2d_cc_w_0_140_s_1_540 = 1.92e-11  mcm5m2d_cf_w_0_140_s_1_540 = 2.31e-11
+ mcm5m2d_ca_w_0_140_s_3_500 = 3.77e-05  mcm5m2d_cc_w_0_140_s_3_500 = 4.21e-12  mcm5m2d_cf_w_0_140_s_3_500 = 3.46e-11
+ mcm5m2d_ca_w_1_120_s_0_140 = 3.77e-05  mcm5m2d_cc_w_1_120_s_0_140 = 1.40e-10  mcm5m2d_cf_w_1_120_s_0_140 = 2.27e-12
+ mcm5m2d_ca_w_1_120_s_0_175 = 3.77e-05  mcm5m2d_cc_w_1_120_s_0_175 = 1.35e-10  mcm5m2d_cf_w_1_120_s_0_175 = 2.93e-12
+ mcm5m2d_ca_w_1_120_s_0_210 = 3.77e-05  mcm5m2d_cc_w_1_120_s_0_210 = 1.27e-10  mcm5m2d_cf_w_1_120_s_0_210 = 3.58e-12
+ mcm5m2d_ca_w_1_120_s_0_280 = 3.77e-05  mcm5m2d_cc_w_1_120_s_0_280 = 1.10e-10  mcm5m2d_cf_w_1_120_s_0_280 = 4.85e-12
+ mcm5m2d_ca_w_1_120_s_0_350 = 3.77e-05  mcm5m2d_cc_w_1_120_s_0_350 = 9.38e-11  mcm5m2d_cf_w_1_120_s_0_350 = 6.12e-12
+ mcm5m2d_ca_w_1_120_s_0_420 = 3.77e-05  mcm5m2d_cc_w_1_120_s_0_420 = 8.12e-11  mcm5m2d_cf_w_1_120_s_0_420 = 7.38e-12
+ mcm5m2d_ca_w_1_120_s_0_560 = 3.77e-05  mcm5m2d_cc_w_1_120_s_0_560 = 6.38e-11  mcm5m2d_cf_w_1_120_s_0_560 = 9.82e-12
+ mcm5m2d_ca_w_1_120_s_0_840 = 3.77e-05  mcm5m2d_cc_w_1_120_s_0_840 = 4.44e-11  mcm5m2d_cf_w_1_120_s_0_840 = 1.44e-11
+ mcm5m2d_ca_w_1_120_s_1_540 = 3.77e-05  mcm5m2d_cc_w_1_120_s_1_540 = 2.28e-11  mcm5m2d_cf_w_1_120_s_1_540 = 2.37e-11
+ mcm5m2d_ca_w_1_120_s_3_500 = 3.77e-05  mcm5m2d_cc_w_1_120_s_3_500 = 5.22e-12  mcm5m2d_cf_w_1_120_s_3_500 = 3.66e-11
+ mcm5m2p1_ca_w_0_140_s_0_140 = 4.39e-05  mcm5m2p1_cc_w_0_140_s_0_140 = 1.18e-10  mcm5m2p1_cf_w_0_140_s_0_140 = 2.59e-12
+ mcm5m2p1_ca_w_0_140_s_0_175 = 4.39e-05  mcm5m2p1_cc_w_0_140_s_0_175 = 1.15e-10  mcm5m2p1_cf_w_0_140_s_0_175 = 3.35e-12
+ mcm5m2p1_ca_w_0_140_s_0_210 = 4.39e-05  mcm5m2p1_cc_w_0_140_s_0_210 = 1.09e-10  mcm5m2p1_cf_w_0_140_s_0_210 = 4.13e-12
+ mcm5m2p1_ca_w_0_140_s_0_280 = 4.39e-05  mcm5m2p1_cc_w_0_140_s_0_280 = 9.36e-11  mcm5m2p1_cf_w_0_140_s_0_280 = 5.63e-12
+ mcm5m2p1_ca_w_0_140_s_0_350 = 4.39e-05  mcm5m2p1_cc_w_0_140_s_0_350 = 7.97e-11  mcm5m2p1_cf_w_0_140_s_0_350 = 7.09e-12
+ mcm5m2p1_ca_w_0_140_s_0_420 = 4.39e-05  mcm5m2p1_cc_w_0_140_s_0_420 = 6.84e-11  mcm5m2p1_cf_w_0_140_s_0_420 = 8.59e-12
+ mcm5m2p1_ca_w_0_140_s_0_560 = 4.39e-05  mcm5m2p1_cc_w_0_140_s_0_560 = 5.32e-11  mcm5m2p1_cf_w_0_140_s_0_560 = 1.14e-11
+ mcm5m2p1_ca_w_0_140_s_0_840 = 4.39e-05  mcm5m2p1_cc_w_0_140_s_0_840 = 3.60e-11  mcm5m2p1_cf_w_0_140_s_0_840 = 1.64e-11
+ mcm5m2p1_ca_w_0_140_s_1_540 = 4.39e-05  mcm5m2p1_cc_w_0_140_s_1_540 = 1.74e-11  mcm5m2p1_cf_w_0_140_s_1_540 = 2.61e-11
+ mcm5m2p1_ca_w_0_140_s_3_500 = 4.39e-05  mcm5m2p1_cc_w_0_140_s_3_500 = 3.36e-12  mcm5m2p1_cf_w_0_140_s_3_500 = 3.74e-11
+ mcm5m2p1_ca_w_1_120_s_0_140 = 4.39e-05  mcm5m2p1_cc_w_1_120_s_0_140 = 1.38e-10  mcm5m2p1_cf_w_1_120_s_0_140 = 2.68e-12
+ mcm5m2p1_ca_w_1_120_s_0_175 = 4.39e-05  mcm5m2p1_cc_w_1_120_s_0_175 = 1.32e-10  mcm5m2p1_cf_w_1_120_s_0_175 = 3.44e-12
+ mcm5m2p1_ca_w_1_120_s_0_210 = 4.39e-05  mcm5m2p1_cc_w_1_120_s_0_210 = 1.24e-10  mcm5m2p1_cf_w_1_120_s_0_210 = 4.20e-12
+ mcm5m2p1_ca_w_1_120_s_0_280 = 4.39e-05  mcm5m2p1_cc_w_1_120_s_0_280 = 1.07e-10  mcm5m2p1_cf_w_1_120_s_0_280 = 5.70e-12
+ mcm5m2p1_ca_w_1_120_s_0_350 = 4.39e-05  mcm5m2p1_cc_w_1_120_s_0_350 = 9.15e-11  mcm5m2p1_cf_w_1_120_s_0_350 = 7.17e-12
+ mcm5m2p1_ca_w_1_120_s_0_420 = 4.39e-05  mcm5m2p1_cc_w_1_120_s_0_420 = 7.92e-11  mcm5m2p1_cf_w_1_120_s_0_420 = 8.62e-12
+ mcm5m2p1_ca_w_1_120_s_0_560 = 4.39e-05  mcm5m2p1_cc_w_1_120_s_0_560 = 6.13e-11  mcm5m2p1_cf_w_1_120_s_0_560 = 1.14e-11
+ mcm5m2p1_ca_w_1_120_s_0_840 = 4.39e-05  mcm5m2p1_cc_w_1_120_s_0_840 = 4.19e-11  mcm5m2p1_cf_w_1_120_s_0_840 = 1.66e-11
+ mcm5m2p1_ca_w_1_120_s_1_540 = 4.39e-05  mcm5m2p1_cc_w_1_120_s_1_540 = 2.06e-11  mcm5m2p1_cf_w_1_120_s_1_540 = 2.67e-11
+ mcm5m2p1_ca_w_1_120_s_3_500 = 4.39e-05  mcm5m2p1_cc_w_1_120_s_3_500 = 4.18e-12  mcm5m2p1_cf_w_1_120_s_3_500 = 3.95e-11
+ mcm5m2l1_ca_w_0_140_s_0_140 = 5.87e-05  mcm5m2l1_cc_w_0_140_s_0_140 = 1.17e-10  mcm5m2l1_cf_w_0_140_s_0_140 = 3.42e-12
+ mcm5m2l1_ca_w_0_140_s_0_175 = 5.87e-05  mcm5m2l1_cc_w_0_140_s_0_175 = 1.13e-10  mcm5m2l1_cf_w_0_140_s_0_175 = 4.44e-12
+ mcm5m2l1_ca_w_0_140_s_0_210 = 5.87e-05  mcm5m2l1_cc_w_0_140_s_0_210 = 1.07e-10  mcm5m2l1_cf_w_0_140_s_0_210 = 5.46e-12
+ mcm5m2l1_ca_w_0_140_s_0_280 = 5.87e-05  mcm5m2l1_cc_w_0_140_s_0_280 = 9.20e-11  mcm5m2l1_cf_w_0_140_s_0_280 = 7.43e-12
+ mcm5m2l1_ca_w_0_140_s_0_350 = 5.87e-05  mcm5m2l1_cc_w_0_140_s_0_350 = 7.72e-11  mcm5m2l1_cf_w_0_140_s_0_350 = 9.36e-12
+ mcm5m2l1_ca_w_0_140_s_0_420 = 5.87e-05  mcm5m2l1_cc_w_0_140_s_0_420 = 6.56e-11  mcm5m2l1_cf_w_0_140_s_0_420 = 1.13e-11
+ mcm5m2l1_ca_w_0_140_s_0_560 = 5.87e-05  mcm5m2l1_cc_w_0_140_s_0_560 = 5.01e-11  mcm5m2l1_cf_w_0_140_s_0_560 = 1.48e-11
+ mcm5m2l1_ca_w_0_140_s_0_840 = 5.87e-05  mcm5m2l1_cc_w_0_140_s_0_840 = 3.27e-11  mcm5m2l1_cf_w_0_140_s_0_840 = 2.11e-11
+ mcm5m2l1_ca_w_0_140_s_1_540 = 5.87e-05  mcm5m2l1_cc_w_0_140_s_1_540 = 1.44e-11  mcm5m2l1_cf_w_0_140_s_1_540 = 3.21e-11
+ mcm5m2l1_ca_w_0_140_s_3_500 = 5.87e-05  mcm5m2l1_cc_w_0_140_s_3_500 = 2.29e-12  mcm5m2l1_cf_w_0_140_s_3_500 = 4.24e-11
+ mcm5m2l1_ca_w_1_120_s_0_140 = 5.87e-05  mcm5m2l1_cc_w_1_120_s_0_140 = 1.35e-10  mcm5m2l1_cf_w_1_120_s_0_140 = 3.46e-12
+ mcm5m2l1_ca_w_1_120_s_0_175 = 5.87e-05  mcm5m2l1_cc_w_1_120_s_0_175 = 1.28e-10  mcm5m2l1_cf_w_1_120_s_0_175 = 4.48e-12
+ mcm5m2l1_ca_w_1_120_s_0_210 = 5.87e-05  mcm5m2l1_cc_w_1_120_s_0_210 = 1.20e-10  mcm5m2l1_cf_w_1_120_s_0_210 = 5.49e-12
+ mcm5m2l1_ca_w_1_120_s_0_280 = 5.87e-05  mcm5m2l1_cc_w_1_120_s_0_280 = 1.03e-10  mcm5m2l1_cf_w_1_120_s_0_280 = 7.47e-12
+ mcm5m2l1_ca_w_1_120_s_0_350 = 5.87e-05  mcm5m2l1_cc_w_1_120_s_0_350 = 8.72e-11  mcm5m2l1_cf_w_1_120_s_0_350 = 9.40e-12
+ mcm5m2l1_ca_w_1_120_s_0_420 = 5.87e-05  mcm5m2l1_cc_w_1_120_s_0_420 = 7.49e-11  mcm5m2l1_cf_w_1_120_s_0_420 = 1.13e-11
+ mcm5m2l1_ca_w_1_120_s_0_560 = 5.87e-05  mcm5m2l1_cc_w_1_120_s_0_560 = 5.72e-11  mcm5m2l1_cf_w_1_120_s_0_560 = 1.49e-11
+ mcm5m2l1_ca_w_1_120_s_0_840 = 5.87e-05  mcm5m2l1_cc_w_1_120_s_0_840 = 3.77e-11  mcm5m2l1_cf_w_1_120_s_0_840 = 2.13e-11
+ mcm5m2l1_ca_w_1_120_s_1_540 = 5.87e-05  mcm5m2l1_cc_w_1_120_s_1_540 = 1.73e-11  mcm5m2l1_cf_w_1_120_s_1_540 = 3.28e-11
+ mcm5m2l1_ca_w_1_120_s_3_500 = 5.87e-05  mcm5m2l1_cc_w_1_120_s_3_500 = 2.99e-12  mcm5m2l1_cf_w_1_120_s_3_500 = 4.48e-11
+ mcm5m2m1_ca_w_0_140_s_0_140 = 2.31e-04  mcm5m2m1_cc_w_0_140_s_0_140 = 1.06e-10  mcm5m2m1_cf_w_0_140_s_0_140 = 1.22e-11
+ mcm5m2m1_ca_w_0_140_s_0_175 = 2.31e-04  mcm5m2m1_cc_w_0_140_s_0_175 = 1.00e-10  mcm5m2m1_cf_w_0_140_s_0_175 = 1.62e-11
+ mcm5m2m1_ca_w_0_140_s_0_210 = 2.31e-04  mcm5m2m1_cc_w_0_140_s_0_210 = 9.28e-11  mcm5m2m1_cf_w_0_140_s_0_210 = 1.99e-11
+ mcm5m2m1_ca_w_0_140_s_0_280 = 2.31e-04  mcm5m2m1_cc_w_0_140_s_0_280 = 7.71e-11  mcm5m2m1_cf_w_0_140_s_0_280 = 2.66e-11
+ mcm5m2m1_ca_w_0_140_s_0_350 = 2.31e-04  mcm5m2m1_cc_w_0_140_s_0_350 = 6.29e-11  mcm5m2m1_cf_w_0_140_s_0_350 = 3.26e-11
+ mcm5m2m1_ca_w_0_140_s_0_420 = 2.31e-04  mcm5m2m1_cc_w_0_140_s_0_420 = 5.12e-11  mcm5m2m1_cf_w_0_140_s_0_420 = 3.78e-11
+ mcm5m2m1_ca_w_0_140_s_0_560 = 2.31e-04  mcm5m2m1_cc_w_0_140_s_0_560 = 3.57e-11  mcm5m2m1_cf_w_0_140_s_0_560 = 4.61e-11
+ mcm5m2m1_ca_w_0_140_s_0_840 = 2.31e-04  mcm5m2m1_cc_w_0_140_s_0_840 = 2.03e-11  mcm5m2m1_cf_w_0_140_s_0_840 = 5.74e-11
+ mcm5m2m1_ca_w_0_140_s_1_540 = 2.31e-04  mcm5m2m1_cc_w_0_140_s_1_540 = 6.76e-12  mcm5m2m1_cf_w_0_140_s_1_540 = 6.98e-11
+ mcm5m2m1_ca_w_0_140_s_3_500 = 2.31e-04  mcm5m2m1_cc_w_0_140_s_3_500 = 7.65e-13  mcm5m2m1_cf_w_0_140_s_3_500 = 7.65e-11
+ mcm5m2m1_ca_w_1_120_s_0_140 = 2.31e-04  mcm5m2m1_cc_w_1_120_s_0_140 = 1.18e-10  mcm5m2m1_cf_w_1_120_s_0_140 = 1.22e-11
+ mcm5m2m1_ca_w_1_120_s_0_175 = 2.31e-04  mcm5m2m1_cc_w_1_120_s_0_175 = 1.11e-10  mcm5m2m1_cf_w_1_120_s_0_175 = 1.62e-11
+ mcm5m2m1_ca_w_1_120_s_0_210 = 2.31e-04  mcm5m2m1_cc_w_1_120_s_0_210 = 1.04e-10  mcm5m2m1_cf_w_1_120_s_0_210 = 1.99e-11
+ mcm5m2m1_ca_w_1_120_s_0_280 = 2.31e-04  mcm5m2m1_cc_w_1_120_s_0_280 = 8.63e-11  mcm5m2m1_cf_w_1_120_s_0_280 = 2.66e-11
+ mcm5m2m1_ca_w_1_120_s_0_350 = 2.31e-04  mcm5m2m1_cc_w_1_120_s_0_350 = 7.07e-11  mcm5m2m1_cf_w_1_120_s_0_350 = 3.25e-11
+ mcm5m2m1_ca_w_1_120_s_0_420 = 2.31e-04  mcm5m2m1_cc_w_1_120_s_0_420 = 5.85e-11  mcm5m2m1_cf_w_1_120_s_0_420 = 3.77e-11
+ mcm5m2m1_ca_w_1_120_s_0_560 = 2.31e-04  mcm5m2m1_cc_w_1_120_s_0_560 = 4.22e-11  mcm5m2m1_cf_w_1_120_s_0_560 = 4.62e-11
+ mcm5m2m1_ca_w_1_120_s_0_840 = 2.31e-04  mcm5m2m1_cc_w_1_120_s_0_840 = 2.50e-11  mcm5m2m1_cf_w_1_120_s_0_840 = 5.77e-11
+ mcm5m2m1_ca_w_1_120_s_1_540 = 2.31e-04  mcm5m2m1_cc_w_1_120_s_1_540 = 9.35e-12  mcm5m2m1_cf_w_1_120_s_1_540 = 7.13e-11
+ mcm5m2m1_ca_w_1_120_s_3_500 = 2.31e-04  mcm5m2m1_cc_w_1_120_s_3_500 = 1.19e-12  mcm5m2m1_cf_w_1_120_s_3_500 = 7.98e-11
+ mcrdlm2f_ca_w_0_140_s_0_140 = 2.53e-05  mcrdlm2f_cc_w_0_140_s_0_140 = 1.22e-10  mcrdlm2f_cf_w_0_140_s_0_140 = 1.50e-12
+ mcrdlm2f_ca_w_0_140_s_0_175 = 2.53e-05  mcrdlm2f_cc_w_0_140_s_0_175 = 1.17e-10  mcrdlm2f_cf_w_0_140_s_0_175 = 1.93e-12
+ mcrdlm2f_ca_w_0_140_s_0_210 = 2.53e-05  mcrdlm2f_cc_w_0_140_s_0_210 = 1.12e-10  mcrdlm2f_cf_w_0_140_s_0_210 = 2.38e-12
+ mcrdlm2f_ca_w_0_140_s_0_280 = 2.53e-05  mcrdlm2f_cc_w_0_140_s_0_280 = 9.65e-11  mcrdlm2f_cf_w_0_140_s_0_280 = 3.25e-12
+ mcrdlm2f_ca_w_0_140_s_0_350 = 2.53e-05  mcrdlm2f_cc_w_0_140_s_0_350 = 8.34e-11  mcrdlm2f_cf_w_0_140_s_0_350 = 4.11e-12
+ mcrdlm2f_ca_w_0_140_s_0_420 = 2.53e-05  mcrdlm2f_cc_w_0_140_s_0_420 = 7.25e-11  mcrdlm2f_cf_w_0_140_s_0_420 = 5.00e-12
+ mcrdlm2f_ca_w_0_140_s_0_560 = 2.53e-05  mcrdlm2f_cc_w_0_140_s_0_560 = 5.79e-11  mcrdlm2f_cf_w_0_140_s_0_560 = 6.63e-12
+ mcrdlm2f_ca_w_0_140_s_0_840 = 2.53e-05  mcrdlm2f_cc_w_0_140_s_0_840 = 4.22e-11  mcrdlm2f_cf_w_0_140_s_0_840 = 9.74e-12
+ mcrdlm2f_ca_w_0_140_s_1_540 = 2.53e-05  mcrdlm2f_cc_w_0_140_s_1_540 = 2.48e-11  mcrdlm2f_cf_w_0_140_s_1_540 = 1.64e-11
+ mcrdlm2f_ca_w_0_140_s_3_500 = 2.53e-05  mcrdlm2f_cc_w_0_140_s_3_500 = 8.90e-12  mcrdlm2f_cf_w_0_140_s_3_500 = 2.72e-11
+ mcrdlm2f_ca_w_1_120_s_0_140 = 2.53e-05  mcrdlm2f_cc_w_1_120_s_0_140 = 1.46e-10  mcrdlm2f_cf_w_1_120_s_0_140 = 1.53e-12
+ mcrdlm2f_ca_w_1_120_s_0_175 = 2.53e-05  mcrdlm2f_cc_w_1_120_s_0_175 = 1.40e-10  mcrdlm2f_cf_w_1_120_s_0_175 = 1.98e-12
+ mcrdlm2f_ca_w_1_120_s_0_210 = 2.53e-05  mcrdlm2f_cc_w_1_120_s_0_210 = 1.33e-10  mcrdlm2f_cf_w_1_120_s_0_210 = 2.42e-12
+ mcrdlm2f_ca_w_1_120_s_0_280 = 2.53e-05  mcrdlm2f_cc_w_1_120_s_0_280 = 1.15e-10  mcrdlm2f_cf_w_1_120_s_0_280 = 3.29e-12
+ mcrdlm2f_ca_w_1_120_s_0_350 = 2.53e-05  mcrdlm2f_cc_w_1_120_s_0_350 = 1.00e-10  mcrdlm2f_cf_w_1_120_s_0_350 = 4.15e-12
+ mcrdlm2f_ca_w_1_120_s_0_420 = 2.53e-05  mcrdlm2f_cc_w_1_120_s_0_420 = 8.84e-11  mcrdlm2f_cf_w_1_120_s_0_420 = 5.00e-12
+ mcrdlm2f_ca_w_1_120_s_0_560 = 2.53e-05  mcrdlm2f_cc_w_1_120_s_0_560 = 7.10e-11  mcrdlm2f_cf_w_1_120_s_0_560 = 6.67e-12
+ mcrdlm2f_ca_w_1_120_s_0_840 = 2.53e-05  mcrdlm2f_cc_w_1_120_s_0_840 = 5.23e-11  mcrdlm2f_cf_w_1_120_s_0_840 = 9.85e-12
+ mcrdlm2f_ca_w_1_120_s_1_540 = 2.53e-05  mcrdlm2f_cc_w_1_120_s_1_540 = 3.14e-11  mcrdlm2f_cf_w_1_120_s_1_540 = 1.68e-11
+ mcrdlm2f_ca_w_1_120_s_3_500 = 2.53e-05  mcrdlm2f_cc_w_1_120_s_3_500 = 1.20e-11  mcrdlm2f_cf_w_1_120_s_3_500 = 2.89e-11
+ mcrdlm2d_ca_w_0_140_s_0_140 = 2.89e-05  mcrdlm2d_cc_w_0_140_s_0_140 = 1.22e-10  mcrdlm2d_cf_w_0_140_s_0_140 = 1.71e-12
+ mcrdlm2d_ca_w_0_140_s_0_175 = 2.89e-05  mcrdlm2d_cc_w_0_140_s_0_175 = 1.17e-10  mcrdlm2d_cf_w_0_140_s_0_175 = 2.21e-12
+ mcrdlm2d_ca_w_0_140_s_0_210 = 2.89e-05  mcrdlm2d_cc_w_0_140_s_0_210 = 1.11e-10  mcrdlm2d_cf_w_0_140_s_0_210 = 2.72e-12
+ mcrdlm2d_ca_w_0_140_s_0_280 = 2.89e-05  mcrdlm2d_cc_w_0_140_s_0_280 = 9.59e-11  mcrdlm2d_cf_w_0_140_s_0_280 = 3.71e-12
+ mcrdlm2d_ca_w_0_140_s_0_350 = 2.89e-05  mcrdlm2d_cc_w_0_140_s_0_350 = 8.27e-11  mcrdlm2d_cf_w_0_140_s_0_350 = 4.69e-12
+ mcrdlm2d_ca_w_0_140_s_0_420 = 2.89e-05  mcrdlm2d_cc_w_0_140_s_0_420 = 7.15e-11  mcrdlm2d_cf_w_0_140_s_0_420 = 5.68e-12
+ mcrdlm2d_ca_w_0_140_s_0_560 = 2.89e-05  mcrdlm2d_cc_w_0_140_s_0_560 = 5.70e-11  mcrdlm2d_cf_w_0_140_s_0_560 = 7.55e-12
+ mcrdlm2d_ca_w_0_140_s_0_840 = 2.89e-05  mcrdlm2d_cc_w_0_140_s_0_840 = 4.10e-11  mcrdlm2d_cf_w_0_140_s_0_840 = 1.10e-11
+ mcrdlm2d_ca_w_0_140_s_1_540 = 2.89e-05  mcrdlm2d_cc_w_0_140_s_1_540 = 2.35e-11  mcrdlm2d_cf_w_0_140_s_1_540 = 1.84e-11
+ mcrdlm2d_ca_w_0_140_s_3_500 = 2.89e-05  mcrdlm2d_cc_w_0_140_s_3_500 = 7.95e-12  mcrdlm2d_cf_w_0_140_s_3_500 = 2.96e-11
+ mcrdlm2d_ca_w_1_120_s_0_140 = 2.89e-05  mcrdlm2d_cc_w_1_120_s_0_140 = 1.44e-10  mcrdlm2d_cf_w_1_120_s_0_140 = 1.76e-12
+ mcrdlm2d_ca_w_1_120_s_0_175 = 2.89e-05  mcrdlm2d_cc_w_1_120_s_0_175 = 1.39e-10  mcrdlm2d_cf_w_1_120_s_0_175 = 2.26e-12
+ mcrdlm2d_ca_w_1_120_s_0_210 = 2.89e-05  mcrdlm2d_cc_w_1_120_s_0_210 = 1.31e-10  mcrdlm2d_cf_w_1_120_s_0_210 = 2.76e-12
+ mcrdlm2d_ca_w_1_120_s_0_280 = 2.89e-05  mcrdlm2d_cc_w_1_120_s_0_280 = 1.13e-10  mcrdlm2d_cf_w_1_120_s_0_280 = 3.75e-12
+ mcrdlm2d_ca_w_1_120_s_0_350 = 2.89e-05  mcrdlm2d_cc_w_1_120_s_0_350 = 9.88e-11  mcrdlm2d_cf_w_1_120_s_0_350 = 4.73e-12
+ mcrdlm2d_ca_w_1_120_s_0_420 = 2.89e-05  mcrdlm2d_cc_w_1_120_s_0_420 = 8.67e-11  mcrdlm2d_cf_w_1_120_s_0_420 = 5.71e-12
+ mcrdlm2d_ca_w_1_120_s_0_560 = 2.89e-05  mcrdlm2d_cc_w_1_120_s_0_560 = 6.94e-11  mcrdlm2d_cf_w_1_120_s_0_560 = 7.59e-12
+ mcrdlm2d_ca_w_1_120_s_0_840 = 2.89e-05  mcrdlm2d_cc_w_1_120_s_0_840 = 5.05e-11  mcrdlm2d_cf_w_1_120_s_0_840 = 1.12e-11
+ mcrdlm2d_ca_w_1_120_s_1_540 = 2.89e-05  mcrdlm2d_cc_w_1_120_s_1_540 = 2.97e-11  mcrdlm2d_cf_w_1_120_s_1_540 = 1.87e-11
+ mcrdlm2d_ca_w_1_120_s_3_500 = 2.89e-05  mcrdlm2d_cc_w_1_120_s_3_500 = 1.08e-11  mcrdlm2d_cf_w_1_120_s_3_500 = 3.14e-11
+ mcrdlm2p1_ca_w_0_140_s_0_140 = 3.52e-05  mcrdlm2p1_cc_w_0_140_s_0_140 = 1.19e-10  mcrdlm2p1_cf_w_0_140_s_0_140 = 2.09e-12
+ mcrdlm2p1_ca_w_0_140_s_0_175 = 3.52e-05  mcrdlm2p1_cc_w_0_140_s_0_175 = 1.16e-10  mcrdlm2p1_cf_w_0_140_s_0_175 = 2.70e-12
+ mcrdlm2p1_ca_w_0_140_s_0_210 = 3.52e-05  mcrdlm2p1_cc_w_0_140_s_0_210 = 1.11e-10  mcrdlm2p1_cf_w_0_140_s_0_210 = 3.31e-12
+ mcrdlm2p1_ca_w_0_140_s_0_280 = 3.52e-05  mcrdlm2p1_cc_w_0_140_s_0_280 = 9.48e-11  mcrdlm2p1_cf_w_0_140_s_0_280 = 4.52e-12
+ mcrdlm2p1_ca_w_0_140_s_0_350 = 3.52e-05  mcrdlm2p1_cc_w_0_140_s_0_350 = 8.16e-11  mcrdlm2p1_cf_w_0_140_s_0_350 = 5.70e-12
+ mcrdlm2p1_ca_w_0_140_s_0_420 = 3.52e-05  mcrdlm2p1_cc_w_0_140_s_0_420 = 7.06e-11  mcrdlm2p1_cf_w_0_140_s_0_420 = 6.90e-12
+ mcrdlm2p1_ca_w_0_140_s_0_560 = 3.52e-05  mcrdlm2p1_cc_w_0_140_s_0_560 = 5.54e-11  mcrdlm2p1_cf_w_0_140_s_0_560 = 9.11e-12
+ mcrdlm2p1_ca_w_0_140_s_0_840 = 3.52e-05  mcrdlm2p1_cc_w_0_140_s_0_840 = 3.93e-11  mcrdlm2p1_cf_w_0_140_s_0_840 = 1.32e-11
+ mcrdlm2p1_ca_w_0_140_s_1_540 = 3.52e-05  mcrdlm2p1_cc_w_0_140_s_1_540 = 2.16e-11  mcrdlm2p1_cf_w_0_140_s_1_540 = 2.15e-11
+ mcrdlm2p1_ca_w_0_140_s_3_500 = 3.52e-05  mcrdlm2p1_cc_w_0_140_s_3_500 = 6.65e-12  mcrdlm2p1_cf_w_0_140_s_3_500 = 3.29e-11
+ mcrdlm2p1_ca_w_1_120_s_0_140 = 3.52e-05  mcrdlm2p1_cc_w_1_120_s_0_140 = 1.42e-10  mcrdlm2p1_cf_w_1_120_s_0_140 = 2.17e-12
+ mcrdlm2p1_ca_w_1_120_s_0_175 = 3.52e-05  mcrdlm2p1_cc_w_1_120_s_0_175 = 1.36e-10  mcrdlm2p1_cf_w_1_120_s_0_175 = 2.79e-12
+ mcrdlm2p1_ca_w_1_120_s_0_210 = 3.52e-05  mcrdlm2p1_cc_w_1_120_s_0_210 = 1.29e-10  mcrdlm2p1_cf_w_1_120_s_0_210 = 3.40e-12
+ mcrdlm2p1_ca_w_1_120_s_0_280 = 3.52e-05  mcrdlm2p1_cc_w_1_120_s_0_280 = 1.11e-10  mcrdlm2p1_cf_w_1_120_s_0_280 = 4.60e-12
+ mcrdlm2p1_ca_w_1_120_s_0_350 = 3.52e-05  mcrdlm2p1_cc_w_1_120_s_0_350 = 9.64e-11  mcrdlm2p1_cf_w_1_120_s_0_350 = 5.78e-12
+ mcrdlm2p1_ca_w_1_120_s_0_420 = 3.52e-05  mcrdlm2p1_cc_w_1_120_s_0_420 = 8.43e-11  mcrdlm2p1_cf_w_1_120_s_0_420 = 6.95e-12
+ mcrdlm2p1_ca_w_1_120_s_0_560 = 3.52e-05  mcrdlm2p1_cc_w_1_120_s_0_560 = 6.70e-11  mcrdlm2p1_cf_w_1_120_s_0_560 = 9.21e-12
+ mcrdlm2p1_ca_w_1_120_s_0_840 = 3.52e-05  mcrdlm2p1_cc_w_1_120_s_0_840 = 4.81e-11  mcrdlm2p1_cf_w_1_120_s_0_840 = 1.34e-11
+ mcrdlm2p1_ca_w_1_120_s_1_540 = 3.52e-05  mcrdlm2p1_cc_w_1_120_s_1_540 = 2.74e-11  mcrdlm2p1_cf_w_1_120_s_1_540 = 2.20e-11
+ mcrdlm2p1_ca_w_1_120_s_3_500 = 3.52e-05  mcrdlm2p1_cc_w_1_120_s_3_500 = 9.37e-12  mcrdlm2p1_cf_w_1_120_s_3_500 = 3.50e-11
+ mcrdlm2l1_ca_w_0_140_s_0_140 = 5.00e-05  mcrdlm2l1_cc_w_0_140_s_0_140 = 1.18e-10  mcrdlm2l1_cf_w_0_140_s_0_140 = 2.91e-12
+ mcrdlm2l1_ca_w_0_140_s_0_175 = 5.00e-05  mcrdlm2l1_cc_w_0_140_s_0_175 = 1.15e-10  mcrdlm2l1_cf_w_0_140_s_0_175 = 3.78e-12
+ mcrdlm2l1_ca_w_0_140_s_0_210 = 5.00e-05  mcrdlm2l1_cc_w_0_140_s_0_210 = 1.08e-10  mcrdlm2l1_cf_w_0_140_s_0_210 = 4.65e-12
+ mcrdlm2l1_ca_w_0_140_s_0_280 = 5.00e-05  mcrdlm2l1_cc_w_0_140_s_0_280 = 9.26e-11  mcrdlm2l1_cf_w_0_140_s_0_280 = 6.33e-12
+ mcrdlm2l1_ca_w_0_140_s_0_350 = 5.00e-05  mcrdlm2l1_cc_w_0_140_s_0_350 = 7.91e-11  mcrdlm2l1_cf_w_0_140_s_0_350 = 7.97e-12
+ mcrdlm2l1_ca_w_0_140_s_0_420 = 5.00e-05  mcrdlm2l1_cc_w_0_140_s_0_420 = 6.78e-11  mcrdlm2l1_cf_w_0_140_s_0_420 = 9.60e-12
+ mcrdlm2l1_ca_w_0_140_s_0_560 = 5.00e-05  mcrdlm2l1_cc_w_0_140_s_0_560 = 5.23e-11  mcrdlm2l1_cf_w_0_140_s_0_560 = 1.26e-11
+ mcrdlm2l1_ca_w_0_140_s_0_840 = 5.00e-05  mcrdlm2l1_cc_w_0_140_s_0_840 = 3.58e-11  mcrdlm2l1_cf_w_0_140_s_0_840 = 1.80e-11
+ mcrdlm2l1_ca_w_0_140_s_1_540 = 5.00e-05  mcrdlm2l1_cc_w_0_140_s_1_540 = 1.82e-11  mcrdlm2l1_cf_w_0_140_s_1_540 = 2.79e-11
+ mcrdlm2l1_ca_w_0_140_s_3_500 = 5.00e-05  mcrdlm2l1_cc_w_0_140_s_3_500 = 4.93e-12  mcrdlm2l1_cf_w_0_140_s_3_500 = 3.91e-11
+ mcrdlm2l1_ca_w_1_120_s_0_140 = 5.00e-05  mcrdlm2l1_cc_w_1_120_s_0_140 = 1.40e-10  mcrdlm2l1_cf_w_1_120_s_0_140 = 2.96e-12
+ mcrdlm2l1_ca_w_1_120_s_0_175 = 5.00e-05  mcrdlm2l1_cc_w_1_120_s_0_175 = 1.32e-10  mcrdlm2l1_cf_w_1_120_s_0_175 = 3.83e-12
+ mcrdlm2l1_ca_w_1_120_s_0_210 = 5.00e-05  mcrdlm2l1_cc_w_1_120_s_0_210 = 1.25e-10  mcrdlm2l1_cf_w_1_120_s_0_210 = 4.69e-12
+ mcrdlm2l1_ca_w_1_120_s_0_280 = 5.00e-05  mcrdlm2l1_cc_w_1_120_s_0_280 = 1.07e-10  mcrdlm2l1_cf_w_1_120_s_0_280 = 6.39e-12
+ mcrdlm2l1_ca_w_1_120_s_0_350 = 5.00e-05  mcrdlm2l1_cc_w_1_120_s_0_350 = 9.25e-11  mcrdlm2l1_cf_w_1_120_s_0_350 = 8.02e-12
+ mcrdlm2l1_ca_w_1_120_s_0_420 = 5.00e-05  mcrdlm2l1_cc_w_1_120_s_0_420 = 8.00e-11  mcrdlm2l1_cf_w_1_120_s_0_420 = 9.62e-12
+ mcrdlm2l1_ca_w_1_120_s_0_560 = 5.00e-05  mcrdlm2l1_cc_w_1_120_s_0_560 = 6.26e-11  mcrdlm2l1_cf_w_1_120_s_0_560 = 1.27e-11
+ mcrdlm2l1_ca_w_1_120_s_0_840 = 5.00e-05  mcrdlm2l1_cc_w_1_120_s_0_840 = 4.40e-11  mcrdlm2l1_cf_w_1_120_s_0_840 = 1.81e-11
+ mcrdlm2l1_ca_w_1_120_s_1_540 = 5.00e-05  mcrdlm2l1_cc_w_1_120_s_1_540 = 2.39e-11  mcrdlm2l1_cf_w_1_120_s_1_540 = 2.85e-11
+ mcrdlm2l1_ca_w_1_120_s_3_500 = 5.00e-05  mcrdlm2l1_cc_w_1_120_s_3_500 = 7.43e-12  mcrdlm2l1_cf_w_1_120_s_3_500 = 4.15e-11
+ mcrdlm2m1_ca_w_0_140_s_0_140 = 2.22e-04  mcrdlm2m1_cc_w_0_140_s_0_140 = 1.07e-10  mcrdlm2m1_cf_w_0_140_s_0_140 = 1.17e-11
+ mcrdlm2m1_ca_w_0_140_s_0_175 = 2.22e-04  mcrdlm2m1_cc_w_0_140_s_0_175 = 1.01e-10  mcrdlm2m1_cf_w_0_140_s_0_175 = 1.55e-11
+ mcrdlm2m1_ca_w_0_140_s_0_210 = 2.22e-04  mcrdlm2m1_cc_w_0_140_s_0_210 = 9.48e-11  mcrdlm2m1_cf_w_0_140_s_0_210 = 1.91e-11
+ mcrdlm2m1_ca_w_0_140_s_0_280 = 2.22e-04  mcrdlm2m1_cc_w_0_140_s_0_280 = 7.84e-11  mcrdlm2m1_cf_w_0_140_s_0_280 = 2.55e-11
+ mcrdlm2m1_ca_w_0_140_s_0_350 = 2.22e-04  mcrdlm2m1_cc_w_0_140_s_0_350 = 6.42e-11  mcrdlm2m1_cf_w_0_140_s_0_350 = 3.11e-11
+ mcrdlm2m1_ca_w_0_140_s_0_420 = 2.22e-04  mcrdlm2m1_cc_w_0_140_s_0_420 = 5.31e-11  mcrdlm2m1_cf_w_0_140_s_0_420 = 3.61e-11
+ mcrdlm2m1_ca_w_0_140_s_0_560 = 2.22e-04  mcrdlm2m1_cc_w_0_140_s_0_560 = 3.81e-11  mcrdlm2m1_cf_w_0_140_s_0_560 = 4.41e-11
+ mcrdlm2m1_ca_w_0_140_s_0_840 = 2.22e-04  mcrdlm2m1_cc_w_0_140_s_0_840 = 2.30e-11  mcrdlm2m1_cf_w_0_140_s_0_840 = 5.47e-11
+ mcrdlm2m1_ca_w_0_140_s_1_540 = 2.22e-04  mcrdlm2m1_cc_w_0_140_s_1_540 = 9.27e-12  mcrdlm2m1_cf_w_0_140_s_1_540 = 6.73e-11
+ mcrdlm2m1_ca_w_0_140_s_3_500 = 2.22e-04  mcrdlm2m1_cc_w_0_140_s_3_500 = 1.97e-12  mcrdlm2m1_cf_w_0_140_s_3_500 = 7.52e-11
+ mcrdlm2m1_ca_w_1_120_s_0_140 = 2.22e-04  mcrdlm2m1_cc_w_1_120_s_0_140 = 1.23e-10  mcrdlm2m1_cf_w_1_120_s_0_140 = 1.17e-11
+ mcrdlm2m1_ca_w_1_120_s_0_175 = 2.22e-04  mcrdlm2m1_cc_w_1_120_s_0_175 = 1.16e-10  mcrdlm2m1_cf_w_1_120_s_0_175 = 1.55e-11
+ mcrdlm2m1_ca_w_1_120_s_0_210 = 2.22e-04  mcrdlm2m1_cc_w_1_120_s_0_210 = 1.08e-10  mcrdlm2m1_cf_w_1_120_s_0_210 = 1.91e-11
+ mcrdlm2m1_ca_w_1_120_s_0_280 = 2.22e-04  mcrdlm2m1_cc_w_1_120_s_0_280 = 9.05e-11  mcrdlm2m1_cf_w_1_120_s_0_280 = 2.56e-11
+ mcrdlm2m1_ca_w_1_120_s_0_350 = 2.22e-04  mcrdlm2m1_cc_w_1_120_s_0_350 = 7.57e-11  mcrdlm2m1_cf_w_1_120_s_0_350 = 3.12e-11
+ mcrdlm2m1_ca_w_1_120_s_0_420 = 2.22e-04  mcrdlm2m1_cc_w_1_120_s_0_420 = 6.41e-11  mcrdlm2m1_cf_w_1_120_s_0_420 = 3.60e-11
+ mcrdlm2m1_ca_w_1_120_s_0_560 = 2.22e-04  mcrdlm2m1_cc_w_1_120_s_0_560 = 4.78e-11  mcrdlm2m1_cf_w_1_120_s_0_560 = 4.41e-11
+ mcrdlm2m1_ca_w_1_120_s_0_840 = 2.22e-04  mcrdlm2m1_cc_w_1_120_s_0_840 = 3.08e-11  mcrdlm2m1_cf_w_1_120_s_0_840 = 5.51e-11
+ mcrdlm2m1_ca_w_1_120_s_1_540 = 2.22e-04  mcrdlm2m1_cc_w_1_120_s_1_540 = 1.46e-11  mcrdlm2m1_cf_w_1_120_s_1_540 = 6.88e-11
+ mcrdlm2m1_ca_w_1_120_s_3_500 = 2.22e-04  mcrdlm2m1_cc_w_1_120_s_3_500 = 3.86e-12  mcrdlm2m1_cf_w_1_120_s_3_500 = 7.94e-11
+ mcm4m3f_ca_w_0_300_s_0_300 = 1.57e-04  mcm4m3f_cc_w_0_300_s_0_300 = 9.81e-11  mcm4m3f_cf_w_0_300_s_0_300 = 1.63e-11
+ mcm4m3f_ca_w_0_300_s_0_360 = 1.57e-04  mcm4m3f_cc_w_0_300_s_0_360 = 8.82e-11  mcm4m3f_cf_w_0_300_s_0_360 = 1.94e-11
+ mcm4m3f_ca_w_0_300_s_0_450 = 1.57e-04  mcm4m3f_cc_w_0_300_s_0_450 = 7.61e-11  mcm4m3f_cf_w_0_300_s_0_450 = 2.37e-11
+ mcm4m3f_ca_w_0_300_s_0_600 = 1.57e-04  mcm4m3f_cc_w_0_300_s_0_600 = 6.02e-11  mcm4m3f_cf_w_0_300_s_0_600 = 2.99e-11
+ mcm4m3f_ca_w_0_300_s_0_800 = 1.57e-04  mcm4m3f_cc_w_0_300_s_0_800 = 4.50e-11  mcm4m3f_cf_w_0_300_s_0_800 = 3.68e-11
+ mcm4m3f_ca_w_0_300_s_1_000 = 1.57e-04  mcm4m3f_cc_w_0_300_s_1_000 = 3.42e-11  mcm4m3f_cf_w_0_300_s_1_000 = 4.26e-11
+ mcm4m3f_ca_w_0_300_s_1_200 = 1.57e-04  mcm4m3f_cc_w_0_300_s_1_200 = 2.64e-11  mcm4m3f_cf_w_0_300_s_1_200 = 4.71e-11
+ mcm4m3f_ca_w_0_300_s_2_100 = 1.57e-04  mcm4m3f_cc_w_0_300_s_2_100 = 9.64e-12  mcm4m3f_cf_w_0_300_s_2_100 = 5.95e-11
+ mcm4m3f_ca_w_0_300_s_3_300 = 1.57e-04  mcm4m3f_cc_w_0_300_s_3_300 = 2.97e-12  mcm4m3f_cf_w_0_300_s_3_300 = 6.56e-11
+ mcm4m3f_ca_w_0_300_s_9_000 = 1.57e-04  mcm4m3f_cc_w_0_300_s_9_000 = 7.00e-14  mcm4m3f_cf_w_0_300_s_9_000 = 6.86e-11
+ mcm4m3f_ca_w_2_400_s_0_300 = 1.57e-04  mcm4m3f_cc_w_2_400_s_0_300 = 1.04e-10  mcm4m3f_cf_w_2_400_s_0_300 = 1.64e-11
+ mcm4m3f_ca_w_2_400_s_0_360 = 1.57e-04  mcm4m3f_cc_w_2_400_s_0_360 = 9.44e-11  mcm4m3f_cf_w_2_400_s_0_360 = 1.95e-11
+ mcm4m3f_ca_w_2_400_s_0_450 = 1.57e-04  mcm4m3f_cc_w_2_400_s_0_450 = 8.13e-11  mcm4m3f_cf_w_2_400_s_0_450 = 2.37e-11
+ mcm4m3f_ca_w_2_400_s_0_600 = 1.57e-04  mcm4m3f_cc_w_2_400_s_0_600 = 6.48e-11  mcm4m3f_cf_w_2_400_s_0_600 = 2.99e-11
+ mcm4m3f_ca_w_2_400_s_0_800 = 1.57e-04  mcm4m3f_cc_w_2_400_s_0_800 = 4.86e-11  mcm4m3f_cf_w_2_400_s_0_800 = 3.69e-11
+ mcm4m3f_ca_w_2_400_s_1_000 = 1.57e-04  mcm4m3f_cc_w_2_400_s_1_000 = 3.70e-11  mcm4m3f_cf_w_2_400_s_1_000 = 4.26e-11
+ mcm4m3f_ca_w_2_400_s_1_200 = 1.57e-04  mcm4m3f_cc_w_2_400_s_1_200 = 2.90e-11  mcm4m3f_cf_w_2_400_s_1_200 = 4.73e-11
+ mcm4m3f_ca_w_2_400_s_2_100 = 1.57e-04  mcm4m3f_cc_w_2_400_s_2_100 = 1.10e-11  mcm4m3f_cf_w_2_400_s_2_100 = 6.02e-11
+ mcm4m3f_ca_w_2_400_s_3_300 = 1.57e-04  mcm4m3f_cc_w_2_400_s_3_300 = 3.52e-12  mcm4m3f_cf_w_2_400_s_3_300 = 6.70e-11
+ mcm4m3f_ca_w_2_400_s_9_000 = 1.57e-04  mcm4m3f_cc_w_2_400_s_9_000 = 3.00e-14  mcm4m3f_cf_w_2_400_s_9_000 = 7.04e-11
+ mcm4m3d_ca_w_0_300_s_0_300 = 1.59e-04  mcm4m3d_cc_w_0_300_s_0_300 = 9.76e-11  mcm4m3d_cf_w_0_300_s_0_300 = 1.65e-11
+ mcm4m3d_ca_w_0_300_s_0_360 = 1.59e-04  mcm4m3d_cc_w_0_300_s_0_360 = 8.78e-11  mcm4m3d_cf_w_0_300_s_0_360 = 1.97e-11
+ mcm4m3d_ca_w_0_300_s_0_450 = 1.59e-04  mcm4m3d_cc_w_0_300_s_0_450 = 7.56e-11  mcm4m3d_cf_w_0_300_s_0_450 = 2.40e-11
+ mcm4m3d_ca_w_0_300_s_0_600 = 1.59e-04  mcm4m3d_cc_w_0_300_s_0_600 = 5.96e-11  mcm4m3d_cf_w_0_300_s_0_600 = 3.04e-11
+ mcm4m3d_ca_w_0_300_s_0_800 = 1.59e-04  mcm4m3d_cc_w_0_300_s_0_800 = 4.44e-11  mcm4m3d_cf_w_0_300_s_0_800 = 3.74e-11
+ mcm4m3d_ca_w_0_300_s_1_000 = 1.59e-04  mcm4m3d_cc_w_0_300_s_1_000 = 3.35e-11  mcm4m3d_cf_w_0_300_s_1_000 = 4.33e-11
+ mcm4m3d_ca_w_0_300_s_1_200 = 1.59e-04  mcm4m3d_cc_w_0_300_s_1_200 = 2.58e-11  mcm4m3d_cf_w_0_300_s_1_200 = 4.79e-11
+ mcm4m3d_ca_w_0_300_s_2_100 = 1.59e-04  mcm4m3d_cc_w_0_300_s_2_100 = 9.03e-12  mcm4m3d_cf_w_0_300_s_2_100 = 6.03e-11
+ mcm4m3d_ca_w_0_300_s_3_300 = 1.59e-04  mcm4m3d_cc_w_0_300_s_3_300 = 2.64e-12  mcm4m3d_cf_w_0_300_s_3_300 = 6.63e-11
+ mcm4m3d_ca_w_0_300_s_9_000 = 1.59e-04  mcm4m3d_cc_w_0_300_s_9_000 = 3.50e-14  mcm4m3d_cf_w_0_300_s_9_000 = 6.89e-11
+ mcm4m3d_ca_w_2_400_s_0_300 = 1.59e-04  mcm4m3d_cc_w_2_400_s_0_300 = 1.03e-10  mcm4m3d_cf_w_2_400_s_0_300 = 1.66e-11
+ mcm4m3d_ca_w_2_400_s_0_360 = 1.59e-04  mcm4m3d_cc_w_2_400_s_0_360 = 9.32e-11  mcm4m3d_cf_w_2_400_s_0_360 = 1.98e-11
+ mcm4m3d_ca_w_2_400_s_0_450 = 1.59e-04  mcm4m3d_cc_w_2_400_s_0_450 = 8.02e-11  mcm4m3d_cf_w_2_400_s_0_450 = 2.41e-11
+ mcm4m3d_ca_w_2_400_s_0_600 = 1.59e-04  mcm4m3d_cc_w_2_400_s_0_600 = 6.37e-11  mcm4m3d_cf_w_2_400_s_0_600 = 3.04e-11
+ mcm4m3d_ca_w_2_400_s_0_800 = 1.59e-04  mcm4m3d_cc_w_2_400_s_0_800 = 4.75e-11  mcm4m3d_cf_w_2_400_s_0_800 = 3.75e-11
+ mcm4m3d_ca_w_2_400_s_1_000 = 1.59e-04  mcm4m3d_cc_w_2_400_s_1_000 = 3.60e-11  mcm4m3d_cf_w_2_400_s_1_000 = 4.34e-11
+ mcm4m3d_ca_w_2_400_s_1_200 = 1.59e-04  mcm4m3d_cc_w_2_400_s_1_200 = 2.78e-11  mcm4m3d_cf_w_2_400_s_1_200 = 4.80e-11
+ mcm4m3d_ca_w_2_400_s_2_100 = 1.59e-04  mcm4m3d_cc_w_2_400_s_2_100 = 1.01e-11  mcm4m3d_cf_w_2_400_s_2_100 = 6.10e-11
+ mcm4m3d_ca_w_2_400_s_3_300 = 1.59e-04  mcm4m3d_cc_w_2_400_s_3_300 = 3.05e-12  mcm4m3d_cf_w_2_400_s_3_300 = 6.75e-11
+ mcm4m3d_ca_w_2_400_s_9_000 = 1.59e-04  mcm4m3d_cc_w_2_400_s_9_000 = 5.50e-14  mcm4m3d_cf_w_2_400_s_9_000 = 7.05e-11
+ mcm4m3p1_ca_w_0_300_s_0_300 = 1.61e-04  mcm4m3p1_cc_w_0_300_s_0_300 = 9.69e-11  mcm4m3p1_cf_w_0_300_s_0_300 = 1.69e-11
+ mcm4m3p1_ca_w_0_300_s_0_360 = 1.61e-04  mcm4m3p1_cc_w_0_300_s_0_360 = 8.71e-11  mcm4m3p1_cf_w_0_300_s_0_360 = 2.01e-11
+ mcm4m3p1_ca_w_0_300_s_0_450 = 1.61e-04  mcm4m3p1_cc_w_0_300_s_0_450 = 7.49e-11  mcm4m3p1_cf_w_0_300_s_0_450 = 2.46e-11
+ mcm4m3p1_ca_w_0_300_s_0_600 = 1.61e-04  mcm4m3p1_cc_w_0_300_s_0_600 = 5.88e-11  mcm4m3p1_cf_w_0_300_s_0_600 = 3.11e-11
+ mcm4m3p1_ca_w_0_300_s_0_800 = 1.61e-04  mcm4m3p1_cc_w_0_300_s_0_800 = 4.35e-11  mcm4m3p1_cf_w_0_300_s_0_800 = 3.83e-11
+ mcm4m3p1_ca_w_0_300_s_1_000 = 1.61e-04  mcm4m3p1_cc_w_0_300_s_1_000 = 3.25e-11  mcm4m3p1_cf_w_0_300_s_1_000 = 4.42e-11
+ mcm4m3p1_ca_w_0_300_s_1_200 = 1.61e-04  mcm4m3p1_cc_w_0_300_s_1_200 = 2.47e-11  mcm4m3p1_cf_w_0_300_s_1_200 = 4.89e-11
+ mcm4m3p1_ca_w_0_300_s_2_100 = 1.61e-04  mcm4m3p1_cc_w_0_300_s_2_100 = 8.20e-12  mcm4m3p1_cf_w_0_300_s_2_100 = 6.15e-11
+ mcm4m3p1_ca_w_0_300_s_3_300 = 1.61e-04  mcm4m3p1_cc_w_0_300_s_3_300 = 2.15e-12  mcm4m3p1_cf_w_0_300_s_3_300 = 6.71e-11
+ mcm4m3p1_ca_w_0_300_s_9_000 = 1.61e-04  mcm4m3p1_cc_w_0_300_s_9_000 = 5.50e-14  mcm4m3p1_cf_w_0_300_s_9_000 = 6.93e-11
+ mcm4m3p1_ca_w_2_400_s_0_300 = 1.61e-04  mcm4m3p1_cc_w_2_400_s_0_300 = 1.02e-10  mcm4m3p1_cf_w_2_400_s_0_300 = 1.70e-11
+ mcm4m3p1_ca_w_2_400_s_0_360 = 1.61e-04  mcm4m3p1_cc_w_2_400_s_0_360 = 9.19e-11  mcm4m3p1_cf_w_2_400_s_0_360 = 2.01e-11
+ mcm4m3p1_ca_w_2_400_s_0_450 = 1.61e-04  mcm4m3p1_cc_w_2_400_s_0_450 = 7.89e-11  mcm4m3p1_cf_w_2_400_s_0_450 = 2.46e-11
+ mcm4m3p1_ca_w_2_400_s_0_600 = 1.61e-04  mcm4m3p1_cc_w_2_400_s_0_600 = 6.21e-11  mcm4m3p1_cf_w_2_400_s_0_600 = 3.11e-11
+ mcm4m3p1_ca_w_2_400_s_0_800 = 1.61e-04  mcm4m3p1_cc_w_2_400_s_0_800 = 4.59e-11  mcm4m3p1_cf_w_2_400_s_0_800 = 3.84e-11
+ mcm4m3p1_ca_w_2_400_s_1_000 = 1.61e-04  mcm4m3p1_cc_w_2_400_s_1_000 = 3.46e-11  mcm4m3p1_cf_w_2_400_s_1_000 = 4.44e-11
+ mcm4m3p1_ca_w_2_400_s_1_200 = 1.61e-04  mcm4m3p1_cc_w_2_400_s_1_200 = 2.63e-11  mcm4m3p1_cf_w_2_400_s_1_200 = 4.92e-11
+ mcm4m3p1_ca_w_2_400_s_2_100 = 1.61e-04  mcm4m3p1_cc_w_2_400_s_2_100 = 8.99e-12  mcm4m3p1_cf_w_2_400_s_2_100 = 6.22e-11
+ mcm4m3p1_ca_w_2_400_s_3_300 = 1.61e-04  mcm4m3p1_cc_w_2_400_s_3_300 = 2.38e-12  mcm4m3p1_cf_w_2_400_s_3_300 = 6.82e-11
+ mcm4m3p1_ca_w_2_400_s_9_000 = 1.61e-04  mcm4m3p1_cc_w_2_400_s_9_000 = 0.00e+00  mcm4m3p1_cf_w_2_400_s_9_000 = 7.07e-11
+ mcm4m3l1_ca_w_0_300_s_0_300 = 1.66e-04  mcm4m3l1_cc_w_0_300_s_0_300 = 9.58e-11  mcm4m3l1_cf_w_0_300_s_0_300 = 1.75e-11
+ mcm4m3l1_ca_w_0_300_s_0_360 = 1.66e-04  mcm4m3l1_cc_w_0_300_s_0_360 = 8.59e-11  mcm4m3l1_cf_w_0_300_s_0_360 = 2.08e-11
+ mcm4m3l1_ca_w_0_300_s_0_450 = 1.66e-04  mcm4m3l1_cc_w_0_300_s_0_450 = 7.36e-11  mcm4m3l1_cf_w_0_300_s_0_450 = 2.54e-11
+ mcm4m3l1_ca_w_0_300_s_0_600 = 1.66e-04  mcm4m3l1_cc_w_0_300_s_0_600 = 5.74e-11  mcm4m3l1_cf_w_0_300_s_0_600 = 3.22e-11
+ mcm4m3l1_ca_w_0_300_s_0_800 = 1.66e-04  mcm4m3l1_cc_w_0_300_s_0_800 = 4.19e-11  mcm4m3l1_cf_w_0_300_s_0_800 = 3.98e-11
+ mcm4m3l1_ca_w_0_300_s_1_000 = 1.66e-04  mcm4m3l1_cc_w_0_300_s_1_000 = 3.09e-11  mcm4m3l1_cf_w_0_300_s_1_000 = 4.60e-11
+ mcm4m3l1_ca_w_0_300_s_1_200 = 1.66e-04  mcm4m3l1_cc_w_0_300_s_1_200 = 2.31e-11  mcm4m3l1_cf_w_0_300_s_1_200 = 5.08e-11
+ mcm4m3l1_ca_w_0_300_s_2_100 = 1.66e-04  mcm4m3l1_cc_w_0_300_s_2_100 = 7.02e-12  mcm4m3l1_cf_w_0_300_s_2_100 = 6.34e-11
+ mcm4m3l1_ca_w_0_300_s_3_300 = 1.66e-04  mcm4m3l1_cc_w_0_300_s_3_300 = 1.64e-12  mcm4m3l1_cf_w_0_300_s_3_300 = 6.85e-11
+ mcm4m3l1_ca_w_0_300_s_9_000 = 1.66e-04  mcm4m3l1_cc_w_0_300_s_9_000 = 1.50e-14  mcm4m3l1_cf_w_0_300_s_9_000 = 7.02e-11
+ mcm4m3l1_ca_w_2_400_s_0_300 = 1.66e-04  mcm4m3l1_cc_w_2_400_s_0_300 = 9.96e-11  mcm4m3l1_cf_w_2_400_s_0_300 = 1.75e-11
+ mcm4m3l1_ca_w_2_400_s_0_360 = 1.66e-04  mcm4m3l1_cc_w_2_400_s_0_360 = 8.95e-11  mcm4m3l1_cf_w_2_400_s_0_360 = 2.08e-11
+ mcm4m3l1_ca_w_2_400_s_0_450 = 1.66e-04  mcm4m3l1_cc_w_2_400_s_0_450 = 7.65e-11  mcm4m3l1_cf_w_2_400_s_0_450 = 2.55e-11
+ mcm4m3l1_ca_w_2_400_s_0_600 = 1.66e-04  mcm4m3l1_cc_w_2_400_s_0_600 = 5.97e-11  mcm4m3l1_cf_w_2_400_s_0_600 = 3.22e-11
+ mcm4m3l1_ca_w_2_400_s_0_800 = 1.66e-04  mcm4m3l1_cc_w_2_400_s_0_800 = 4.37e-11  mcm4m3l1_cf_w_2_400_s_0_800 = 3.99e-11
+ mcm4m3l1_ca_w_2_400_s_1_000 = 1.66e-04  mcm4m3l1_cc_w_2_400_s_1_000 = 3.23e-11  mcm4m3l1_cf_w_2_400_s_1_000 = 4.61e-11
+ mcm4m3l1_ca_w_2_400_s_1_200 = 1.66e-04  mcm4m3l1_cc_w_2_400_s_1_200 = 2.42e-11  mcm4m3l1_cf_w_2_400_s_1_200 = 5.11e-11
+ mcm4m3l1_ca_w_2_400_s_2_100 = 1.66e-04  mcm4m3l1_cc_w_2_400_s_2_100 = 7.42e-12  mcm4m3l1_cf_w_2_400_s_2_100 = 6.40e-11
+ mcm4m3l1_ca_w_2_400_s_3_300 = 1.66e-04  mcm4m3l1_cc_w_2_400_s_3_300 = 1.74e-12  mcm4m3l1_cf_w_2_400_s_3_300 = 6.94e-11
+ mcm4m3l1_ca_w_2_400_s_9_000 = 1.66e-04  mcm4m3l1_cc_w_2_400_s_9_000 = 2.00e-14  mcm4m3l1_cf_w_2_400_s_9_000 = 7.12e-11
+ mcm4m3m1_ca_w_0_300_s_0_300 = 1.83e-04  mcm4m3m1_cc_w_0_300_s_0_300 = 9.22e-11  mcm4m3m1_cf_w_0_300_s_0_300 = 1.95e-11
+ mcm4m3m1_ca_w_0_300_s_0_360 = 1.83e-04  mcm4m3m1_cc_w_0_300_s_0_360 = 8.23e-11  mcm4m3m1_cf_w_0_300_s_0_360 = 2.33e-11
+ mcm4m3m1_ca_w_0_300_s_0_450 = 1.83e-04  mcm4m3m1_cc_w_0_300_s_0_450 = 6.96e-11  mcm4m3m1_cf_w_0_300_s_0_450 = 2.85e-11
+ mcm4m3m1_ca_w_0_300_s_0_600 = 1.83e-04  mcm4m3m1_cc_w_0_300_s_0_600 = 5.32e-11  mcm4m3m1_cf_w_0_300_s_0_600 = 3.62e-11
+ mcm4m3m1_ca_w_0_300_s_0_800 = 1.83e-04  mcm4m3m1_cc_w_0_300_s_0_800 = 3.75e-11  mcm4m3m1_cf_w_0_300_s_0_800 = 4.47e-11
+ mcm4m3m1_ca_w_0_300_s_1_000 = 1.83e-04  mcm4m3m1_cc_w_0_300_s_1_000 = 2.64e-11  mcm4m3m1_cf_w_0_300_s_1_000 = 5.16e-11
+ mcm4m3m1_ca_w_0_300_s_1_200 = 1.83e-04  mcm4m3m1_cc_w_0_300_s_1_200 = 1.88e-11  mcm4m3m1_cf_w_0_300_s_1_200 = 5.69e-11
+ mcm4m3m1_ca_w_0_300_s_2_100 = 1.83e-04  mcm4m3m1_cc_w_0_300_s_2_100 = 4.46e-12  mcm4m3m1_cf_w_0_300_s_2_100 = 6.91e-11
+ mcm4m3m1_ca_w_0_300_s_3_300 = 1.83e-04  mcm4m3m1_cc_w_0_300_s_3_300 = 7.10e-13  mcm4m3m1_cf_w_0_300_s_3_300 = 7.28e-11
+ mcm4m3m1_ca_w_0_300_s_9_000 = 1.83e-04  mcm4m3m1_cc_w_0_300_s_9_000 = 6.00e-14  mcm4m3m1_cf_w_0_300_s_9_000 = 7.35e-11
+ mcm4m3m1_ca_w_2_400_s_0_300 = 1.83e-04  mcm4m3m1_cc_w_2_400_s_0_300 = 9.36e-11  mcm4m3m1_cf_w_2_400_s_0_300 = 1.96e-11
+ mcm4m3m1_ca_w_2_400_s_0_360 = 1.83e-04  mcm4m3m1_cc_w_2_400_s_0_360 = 8.36e-11  mcm4m3m1_cf_w_2_400_s_0_360 = 2.33e-11
+ mcm4m3m1_ca_w_2_400_s_0_450 = 1.83e-04  mcm4m3m1_cc_w_2_400_s_0_450 = 7.08e-11  mcm4m3m1_cf_w_2_400_s_0_450 = 2.85e-11
+ mcm4m3m1_ca_w_2_400_s_0_600 = 1.83e-04  mcm4m3m1_cc_w_2_400_s_0_600 = 5.41e-11  mcm4m3m1_cf_w_2_400_s_0_600 = 3.62e-11
+ mcm4m3m1_ca_w_2_400_s_0_800 = 1.83e-04  mcm4m3m1_cc_w_2_400_s_0_800 = 3.81e-11  mcm4m3m1_cf_w_2_400_s_0_800 = 4.48e-11
+ mcm4m3m1_ca_w_2_400_s_1_000 = 1.83e-04  mcm4m3m1_cc_w_2_400_s_1_000 = 2.69e-11  mcm4m3m1_cf_w_2_400_s_1_000 = 5.17e-11
+ mcm4m3m1_ca_w_2_400_s_1_200 = 1.83e-04  mcm4m3m1_cc_w_2_400_s_1_200 = 1.92e-11  mcm4m3m1_cf_w_2_400_s_1_200 = 5.70e-11
+ mcm4m3m1_ca_w_2_400_s_2_100 = 1.83e-04  mcm4m3m1_cc_w_2_400_s_2_100 = 4.55e-12  mcm4m3m1_cf_w_2_400_s_2_100 = 6.93e-11
+ mcm4m3m1_ca_w_2_400_s_3_300 = 1.83e-04  mcm4m3m1_cc_w_2_400_s_3_300 = 7.50e-13  mcm4m3m1_cf_w_2_400_s_3_300 = 7.31e-11
+ mcm4m3m1_ca_w_2_400_s_9_000 = 1.83e-04  mcm4m3m1_cc_w_2_400_s_9_000 = 0.00e+00  mcm4m3m1_cf_w_2_400_s_9_000 = 7.39e-11
+ mcm4m3m2_ca_w_0_300_s_0_300 = 2.54e-04  mcm4m3m2_cc_w_0_300_s_0_300 = 8.27e-11  mcm4m3m2_cf_w_0_300_s_0_300 = 2.75e-11
+ mcm4m3m2_ca_w_0_300_s_0_360 = 2.54e-04  mcm4m3m2_cc_w_0_300_s_0_360 = 7.25e-11  mcm4m3m2_cf_w_0_300_s_0_360 = 3.27e-11
+ mcm4m3m2_ca_w_0_300_s_0_450 = 2.54e-04  mcm4m3m2_cc_w_0_300_s_0_450 = 6.00e-11  mcm4m3m2_cf_w_0_300_s_0_450 = 3.98e-11
+ mcm4m3m2_ca_w_0_300_s_0_600 = 2.54e-04  mcm4m3m2_cc_w_0_300_s_0_600 = 4.36e-11  mcm4m3m2_cf_w_0_300_s_0_600 = 4.98e-11
+ mcm4m3m2_ca_w_0_300_s_0_800 = 2.54e-04  mcm4m3m2_cc_w_0_300_s_0_800 = 2.87e-11  mcm4m3m2_cf_w_0_300_s_0_800 = 6.04e-11
+ mcm4m3m2_ca_w_0_300_s_1_000 = 2.54e-04  mcm4m3m2_cc_w_0_300_s_1_000 = 1.85e-11  mcm4m3m2_cf_w_0_300_s_1_000 = 6.87e-11
+ mcm4m3m2_ca_w_0_300_s_1_200 = 2.54e-04  mcm4m3m2_cc_w_0_300_s_1_200 = 1.19e-11  mcm4m3m2_cf_w_0_300_s_1_200 = 7.38e-11
+ mcm4m3m2_ca_w_0_300_s_2_100 = 2.54e-04  mcm4m3m2_cc_w_0_300_s_2_100 = 1.80e-12  mcm4m3m2_cf_w_0_300_s_2_100 = 8.36e-11
+ mcm4m3m2_ca_w_0_300_s_3_300 = 2.54e-04  mcm4m3m2_cc_w_0_300_s_3_300 = 2.00e-13  mcm4m3m2_cf_w_0_300_s_3_300 = 8.52e-11
+ mcm4m3m2_ca_w_0_300_s_9_000 = 2.54e-04  mcm4m3m2_cc_w_0_300_s_9_000 = 0.00e+00  mcm4m3m2_cf_w_0_300_s_9_000 = 8.54e-11
+ mcm4m3m2_ca_w_2_400_s_0_300 = 2.54e-04  mcm4m3m2_cc_w_2_400_s_0_300 = 8.29e-11  mcm4m3m2_cf_w_2_400_s_0_300 = 2.75e-11
+ mcm4m3m2_ca_w_2_400_s_0_360 = 2.54e-04  mcm4m3m2_cc_w_2_400_s_0_360 = 7.29e-11  mcm4m3m2_cf_w_2_400_s_0_360 = 3.27e-11
+ mcm4m3m2_ca_w_2_400_s_0_450 = 2.54e-04  mcm4m3m2_cc_w_2_400_s_0_450 = 6.03e-11  mcm4m3m2_cf_w_2_400_s_0_450 = 3.98e-11
+ mcm4m3m2_ca_w_2_400_s_0_600 = 2.54e-04  mcm4m3m2_cc_w_2_400_s_0_600 = 4.40e-11  mcm4m3m2_cf_w_2_400_s_0_600 = 4.99e-11
+ mcm4m3m2_ca_w_2_400_s_0_800 = 2.54e-04  mcm4m3m2_cc_w_2_400_s_0_800 = 2.88e-11  mcm4m3m2_cf_w_2_400_s_0_800 = 6.05e-11
+ mcm4m3m2_ca_w_2_400_s_1_000 = 2.54e-04  mcm4m3m2_cc_w_2_400_s_1_000 = 1.86e-11  mcm4m3m2_cf_w_2_400_s_1_000 = 6.85e-11
+ mcm4m3m2_ca_w_2_400_s_1_200 = 2.54e-04  mcm4m3m2_cc_w_2_400_s_1_200 = 1.19e-11  mcm4m3m2_cf_w_2_400_s_1_200 = 7.40e-11
+ mcm4m3m2_ca_w_2_400_s_2_100 = 2.54e-04  mcm4m3m2_cc_w_2_400_s_2_100 = 1.75e-12  mcm4m3m2_cf_w_2_400_s_2_100 = 8.36e-11
+ mcm4m3m2_ca_w_2_400_s_3_300 = 2.54e-04  mcm4m3m2_cc_w_2_400_s_3_300 = 2.00e-13  mcm4m3m2_cf_w_2_400_s_3_300 = 8.55e-11
+ mcm4m3m2_ca_w_2_400_s_9_000 = 2.54e-04  mcm4m3m2_cc_w_2_400_s_9_000 = 0.00e+00  mcm4m3m2_cf_w_2_400_s_9_000 = 8.57e-11
+ mcm5m3f_ca_w_0_300_s_0_300 = 3.79e-05  mcm5m3f_cc_w_0_300_s_0_300 = 1.13e-10  mcm5m3f_cf_w_0_300_s_0_300 = 4.89e-12
+ mcm5m3f_ca_w_0_300_s_0_360 = 3.79e-05  mcm5m3f_cc_w_0_300_s_0_360 = 1.04e-10  mcm5m3f_cf_w_0_300_s_0_360 = 5.97e-12
+ mcm5m3f_ca_w_0_300_s_0_450 = 3.79e-05  mcm5m3f_cc_w_0_300_s_0_450 = 9.13e-11  mcm5m3f_cf_w_0_300_s_0_450 = 7.59e-12
+ mcm5m3f_ca_w_0_300_s_0_600 = 3.79e-05  mcm5m3f_cc_w_0_300_s_0_600 = 7.55e-11  mcm5m3f_cf_w_0_300_s_0_600 = 1.02e-11
+ mcm5m3f_ca_w_0_300_s_0_800 = 3.79e-05  mcm5m3f_cc_w_0_300_s_0_800 = 6.00e-11  mcm5m3f_cf_w_0_300_s_0_800 = 1.34e-11
+ mcm5m3f_ca_w_0_300_s_1_000 = 3.79e-05  mcm5m3f_cc_w_0_300_s_1_000 = 4.86e-11  mcm5m3f_cf_w_0_300_s_1_000 = 1.65e-11
+ mcm5m3f_ca_w_0_300_s_1_200 = 3.79e-05  mcm5m3f_cc_w_0_300_s_1_200 = 4.01e-11  mcm5m3f_cf_w_0_300_s_1_200 = 1.94e-11
+ mcm5m3f_ca_w_0_300_s_2_100 = 3.79e-05  mcm5m3f_cc_w_0_300_s_2_100 = 1.95e-11  mcm5m3f_cf_w_0_300_s_2_100 = 2.99e-11
+ mcm5m3f_ca_w_0_300_s_3_300 = 3.79e-05  mcm5m3f_cc_w_0_300_s_3_300 = 8.30e-12  mcm5m3f_cf_w_0_300_s_3_300 = 3.81e-11
+ mcm5m3f_ca_w_0_300_s_9_000 = 3.79e-05  mcm5m3f_cc_w_0_300_s_9_000 = 2.00e-13  mcm5m3f_cf_w_0_300_s_9_000 = 4.56e-11
+ mcm5m3f_ca_w_2_400_s_0_300 = 3.79e-05  mcm5m3f_cc_w_2_400_s_0_300 = 1.23e-10  mcm5m3f_cf_w_2_400_s_0_300 = 4.95e-12
+ mcm5m3f_ca_w_2_400_s_0_360 = 3.79e-05  mcm5m3f_cc_w_2_400_s_0_360 = 1.13e-10  mcm5m3f_cf_w_2_400_s_0_360 = 6.01e-12
+ mcm5m3f_ca_w_2_400_s_0_450 = 3.79e-05  mcm5m3f_cc_w_2_400_s_0_450 = 1.00e-10  mcm5m3f_cf_w_2_400_s_0_450 = 7.61e-12
+ mcm5m3f_ca_w_2_400_s_0_600 = 3.79e-05  mcm5m3f_cc_w_2_400_s_0_600 = 8.25e-11  mcm5m3f_cf_w_2_400_s_0_600 = 1.02e-11
+ mcm5m3f_ca_w_2_400_s_0_800 = 3.79e-05  mcm5m3f_cc_w_2_400_s_0_800 = 6.56e-11  mcm5m3f_cf_w_2_400_s_0_800 = 1.35e-11
+ mcm5m3f_ca_w_2_400_s_1_000 = 3.79e-05  mcm5m3f_cc_w_2_400_s_1_000 = 5.31e-11  mcm5m3f_cf_w_2_400_s_1_000 = 1.67e-11
+ mcm5m3f_ca_w_2_400_s_1_200 = 3.79e-05  mcm5m3f_cc_w_2_400_s_1_200 = 4.38e-11  mcm5m3f_cf_w_2_400_s_1_200 = 1.96e-11
+ mcm5m3f_ca_w_2_400_s_2_100 = 3.79e-05  mcm5m3f_cc_w_2_400_s_2_100 = 2.14e-11  mcm5m3f_cf_w_2_400_s_2_100 = 3.05e-11
+ mcm5m3f_ca_w_2_400_s_3_300 = 3.79e-05  mcm5m3f_cc_w_2_400_s_3_300 = 9.27e-12  mcm5m3f_cf_w_2_400_s_3_300 = 3.93e-11
+ mcm5m3f_ca_w_2_400_s_9_000 = 3.79e-05  mcm5m3f_cc_w_2_400_s_9_000 = 2.55e-13  mcm5m3f_cf_w_2_400_s_9_000 = 4.77e-11
+ mcm5m3d_ca_w_0_300_s_0_300 = 3.96e-05  mcm5m3d_cc_w_0_300_s_0_300 = 1.13e-10  mcm5m3d_cf_w_0_300_s_0_300 = 5.12e-12
+ mcm5m3d_ca_w_0_300_s_0_360 = 3.96e-05  mcm5m3d_cc_w_0_300_s_0_360 = 1.03e-10  mcm5m3d_cf_w_0_300_s_0_360 = 6.24e-12
+ mcm5m3d_ca_w_0_300_s_0_450 = 3.96e-05  mcm5m3d_cc_w_0_300_s_0_450 = 9.08e-11  mcm5m3d_cf_w_0_300_s_0_450 = 7.93e-12
+ mcm5m3d_ca_w_0_300_s_0_600 = 3.96e-05  mcm5m3d_cc_w_0_300_s_0_600 = 7.50e-11  mcm5m3d_cf_w_0_300_s_0_600 = 1.06e-11
+ mcm5m3d_ca_w_0_300_s_0_800 = 3.96e-05  mcm5m3d_cc_w_0_300_s_0_800 = 5.94e-11  mcm5m3d_cf_w_0_300_s_0_800 = 1.40e-11
+ mcm5m3d_ca_w_0_300_s_1_000 = 3.96e-05  mcm5m3d_cc_w_0_300_s_1_000 = 4.79e-11  mcm5m3d_cf_w_0_300_s_1_000 = 1.72e-11
+ mcm5m3d_ca_w_0_300_s_1_200 = 3.96e-05  mcm5m3d_cc_w_0_300_s_1_200 = 3.93e-11  mcm5m3d_cf_w_0_300_s_1_200 = 2.02e-11
+ mcm5m3d_ca_w_0_300_s_2_100 = 3.96e-05  mcm5m3d_cc_w_0_300_s_2_100 = 1.87e-11  mcm5m3d_cf_w_0_300_s_2_100 = 3.10e-11
+ mcm5m3d_ca_w_0_300_s_3_300 = 3.96e-05  mcm5m3d_cc_w_0_300_s_3_300 = 7.73e-12  mcm5m3d_cf_w_0_300_s_3_300 = 3.93e-11
+ mcm5m3d_ca_w_0_300_s_9_000 = 3.96e-05  mcm5m3d_cc_w_0_300_s_9_000 = 1.75e-13  mcm5m3d_cf_w_0_300_s_9_000 = 4.62e-11
+ mcm5m3d_ca_w_2_400_s_0_300 = 3.96e-05  mcm5m3d_cc_w_2_400_s_0_300 = 1.22e-10  mcm5m3d_cf_w_2_400_s_0_300 = 5.17e-12
+ mcm5m3d_ca_w_2_400_s_0_360 = 3.96e-05  mcm5m3d_cc_w_2_400_s_0_360 = 1.12e-10  mcm5m3d_cf_w_2_400_s_0_360 = 6.29e-12
+ mcm5m3d_ca_w_2_400_s_0_450 = 3.96e-05  mcm5m3d_cc_w_2_400_s_0_450 = 9.88e-11  mcm5m3d_cf_w_2_400_s_0_450 = 7.95e-12
+ mcm5m3d_ca_w_2_400_s_0_600 = 3.96e-05  mcm5m3d_cc_w_2_400_s_0_600 = 8.13e-11  mcm5m3d_cf_w_2_400_s_0_600 = 1.07e-11
+ mcm5m3d_ca_w_2_400_s_0_800 = 3.96e-05  mcm5m3d_cc_w_2_400_s_0_800 = 6.44e-11  mcm5m3d_cf_w_2_400_s_0_800 = 1.41e-11
+ mcm5m3d_ca_w_2_400_s_1_000 = 3.96e-05  mcm5m3d_cc_w_2_400_s_1_000 = 5.20e-11  mcm5m3d_cf_w_2_400_s_1_000 = 1.74e-11
+ mcm5m3d_ca_w_2_400_s_1_200 = 3.96e-05  mcm5m3d_cc_w_2_400_s_1_200 = 4.27e-11  mcm5m3d_cf_w_2_400_s_1_200 = 2.05e-11
+ mcm5m3d_ca_w_2_400_s_2_100 = 3.96e-05  mcm5m3d_cc_w_2_400_s_2_100 = 2.04e-11  mcm5m3d_cf_w_2_400_s_2_100 = 3.16e-11
+ mcm5m3d_ca_w_2_400_s_3_300 = 3.96e-05  mcm5m3d_cc_w_2_400_s_3_300 = 8.54e-12  mcm5m3d_cf_w_2_400_s_3_300 = 4.04e-11
+ mcm5m3d_ca_w_2_400_s_9_000 = 3.96e-05  mcm5m3d_cc_w_2_400_s_9_000 = 1.75e-13  mcm5m3d_cf_w_2_400_s_9_000 = 4.81e-11
+ mcm5m3p1_ca_w_0_300_s_0_300 = 4.22e-05  mcm5m3p1_cc_w_0_300_s_0_300 = 1.12e-10  mcm5m3p1_cf_w_0_300_s_0_300 = 5.46e-12
+ mcm5m3p1_ca_w_0_300_s_0_360 = 4.22e-05  mcm5m3p1_cc_w_0_300_s_0_360 = 1.02e-10  mcm5m3p1_cf_w_0_300_s_0_360 = 6.66e-12
+ mcm5m3p1_ca_w_0_300_s_0_450 = 4.22e-05  mcm5m3p1_cc_w_0_300_s_0_450 = 9.01e-11  mcm5m3p1_cf_w_0_300_s_0_450 = 8.44e-12
+ mcm5m3p1_ca_w_0_300_s_0_600 = 4.22e-05  mcm5m3p1_cc_w_0_300_s_0_600 = 7.41e-11  mcm5m3p1_cf_w_0_300_s_0_600 = 1.13e-11
+ mcm5m3p1_ca_w_0_300_s_0_800 = 4.22e-05  mcm5m3p1_cc_w_0_300_s_0_800 = 5.84e-11  mcm5m3p1_cf_w_0_300_s_0_800 = 1.49e-11
+ mcm5m3p1_ca_w_0_300_s_1_000 = 4.22e-05  mcm5m3p1_cc_w_0_300_s_1_000 = 4.69e-11  mcm5m3p1_cf_w_0_300_s_1_000 = 1.83e-11
+ mcm5m3p1_ca_w_0_300_s_1_200 = 4.22e-05  mcm5m3p1_cc_w_0_300_s_1_200 = 3.83e-11  mcm5m3p1_cf_w_0_300_s_1_200 = 2.15e-11
+ mcm5m3p1_ca_w_0_300_s_2_100 = 4.22e-05  mcm5m3p1_cc_w_0_300_s_2_100 = 1.75e-11  mcm5m3p1_cf_w_0_300_s_2_100 = 3.26e-11
+ mcm5m3p1_ca_w_0_300_s_3_300 = 4.22e-05  mcm5m3p1_cc_w_0_300_s_3_300 = 6.94e-12  mcm5m3p1_cf_w_0_300_s_3_300 = 4.09e-11
+ mcm5m3p1_ca_w_0_300_s_9_000 = 4.22e-05  mcm5m3p1_cc_w_0_300_s_9_000 = 1.25e-13  mcm5m3p1_cf_w_0_300_s_9_000 = 4.72e-11
+ mcm5m3p1_ca_w_2_400_s_0_300 = 4.22e-05  mcm5m3p1_cc_w_2_400_s_0_300 = 1.21e-10  mcm5m3p1_cf_w_2_400_s_0_300 = 5.55e-12
+ mcm5m3p1_ca_w_2_400_s_0_360 = 4.22e-05  mcm5m3p1_cc_w_2_400_s_0_360 = 1.11e-10  mcm5m3p1_cf_w_2_400_s_0_360 = 6.74e-12
+ mcm5m3p1_ca_w_2_400_s_0_450 = 4.22e-05  mcm5m3p1_cc_w_2_400_s_0_450 = 9.73e-11  mcm5m3p1_cf_w_2_400_s_0_450 = 8.51e-12
+ mcm5m3p1_ca_w_2_400_s_0_600 = 4.22e-05  mcm5m3p1_cc_w_2_400_s_0_600 = 7.98e-11  mcm5m3p1_cf_w_2_400_s_0_600 = 1.14e-11
+ mcm5m3p1_ca_w_2_400_s_0_800 = 4.22e-05  mcm5m3p1_cc_w_2_400_s_0_800 = 6.29e-11  mcm5m3p1_cf_w_2_400_s_0_800 = 1.50e-11
+ mcm5m3p1_ca_w_2_400_s_1_000 = 4.22e-05  mcm5m3p1_cc_w_2_400_s_1_000 = 5.04e-11  mcm5m3p1_cf_w_2_400_s_1_000 = 1.85e-11
+ mcm5m3p1_ca_w_2_400_s_1_200 = 4.22e-05  mcm5m3p1_cc_w_2_400_s_1_200 = 4.11e-11  mcm5m3p1_cf_w_2_400_s_1_200 = 2.18e-11
+ mcm5m3p1_ca_w_2_400_s_2_100 = 4.22e-05  mcm5m3p1_cc_w_2_400_s_2_100 = 1.90e-11  mcm5m3p1_cf_w_2_400_s_2_100 = 3.33e-11
+ mcm5m3p1_ca_w_2_400_s_3_300 = 4.22e-05  mcm5m3p1_cc_w_2_400_s_3_300 = 7.50e-12  mcm5m3p1_cf_w_2_400_s_3_300 = 4.20e-11
+ mcm5m3p1_ca_w_2_400_s_9_000 = 4.22e-05  mcm5m3p1_cc_w_2_400_s_9_000 = 1.25e-13  mcm5m3p1_cf_w_2_400_s_9_000 = 4.89e-11
+ mcm5m3l1_ca_w_0_300_s_0_300 = 4.70e-05  mcm5m3l1_cc_w_0_300_s_0_300 = 1.11e-10  mcm5m3l1_cf_w_0_300_s_0_300 = 6.05e-12
+ mcm5m3l1_ca_w_0_300_s_0_360 = 4.70e-05  mcm5m3l1_cc_w_0_300_s_0_360 = 1.01e-10  mcm5m3l1_cf_w_0_300_s_0_360 = 7.37e-12
+ mcm5m3l1_ca_w_0_300_s_0_450 = 4.70e-05  mcm5m3l1_cc_w_0_300_s_0_450 = 8.88e-11  mcm5m3l1_cf_w_0_300_s_0_450 = 9.33e-12
+ mcm5m3l1_ca_w_0_300_s_0_600 = 4.70e-05  mcm5m3l1_cc_w_0_300_s_0_600 = 7.27e-11  mcm5m3l1_cf_w_0_300_s_0_600 = 1.25e-11
+ mcm5m3l1_ca_w_0_300_s_0_800 = 4.70e-05  mcm5m3l1_cc_w_0_300_s_0_800 = 5.69e-11  mcm5m3l1_cf_w_0_300_s_0_800 = 1.64e-11
+ mcm5m3l1_ca_w_0_300_s_1_000 = 4.70e-05  mcm5m3l1_cc_w_0_300_s_1_000 = 4.52e-11  mcm5m3l1_cf_w_0_300_s_1_000 = 2.02e-11
+ mcm5m3l1_ca_w_0_300_s_1_200 = 4.70e-05  mcm5m3l1_cc_w_0_300_s_1_200 = 3.66e-11  mcm5m3l1_cf_w_0_300_s_1_200 = 2.35e-11
+ mcm5m3l1_ca_w_0_300_s_2_100 = 4.70e-05  mcm5m3l1_cc_w_0_300_s_2_100 = 1.59e-11  mcm5m3l1_cf_w_0_300_s_2_100 = 3.52e-11
+ mcm5m3l1_ca_w_0_300_s_3_300 = 4.70e-05  mcm5m3l1_cc_w_0_300_s_3_300 = 5.83e-12  mcm5m3l1_cf_w_0_300_s_3_300 = 4.34e-11
+ mcm5m3l1_ca_w_0_300_s_9_000 = 4.70e-05  mcm5m3l1_cc_w_0_300_s_9_000 = 1.10e-13  mcm5m3l1_cf_w_0_300_s_9_000 = 4.89e-11
+ mcm5m3l1_ca_w_2_400_s_0_300 = 4.70e-05  mcm5m3l1_cc_w_2_400_s_0_300 = 1.19e-10  mcm5m3l1_cf_w_2_400_s_0_300 = 6.09e-12
+ mcm5m3l1_ca_w_2_400_s_0_360 = 4.70e-05  mcm5m3l1_cc_w_2_400_s_0_360 = 1.08e-10  mcm5m3l1_cf_w_2_400_s_0_360 = 7.41e-12
+ mcm5m3l1_ca_w_2_400_s_0_450 = 4.70e-05  mcm5m3l1_cc_w_2_400_s_0_450 = 9.46e-11  mcm5m3l1_cf_w_2_400_s_0_450 = 9.36e-12
+ mcm5m3l1_ca_w_2_400_s_0_600 = 4.70e-05  mcm5m3l1_cc_w_2_400_s_0_600 = 7.73e-11  mcm5m3l1_cf_w_2_400_s_0_600 = 1.25e-11
+ mcm5m3l1_ca_w_2_400_s_0_800 = 4.70e-05  mcm5m3l1_cc_w_2_400_s_0_800 = 6.06e-11  mcm5m3l1_cf_w_2_400_s_0_800 = 1.65e-11
+ mcm5m3l1_ca_w_2_400_s_1_000 = 4.70e-05  mcm5m3l1_cc_w_2_400_s_1_000 = 4.81e-11  mcm5m3l1_cf_w_2_400_s_1_000 = 2.04e-11
+ mcm5m3l1_ca_w_2_400_s_1_200 = 4.70e-05  mcm5m3l1_cc_w_2_400_s_1_200 = 3.89e-11  mcm5m3l1_cf_w_2_400_s_1_200 = 2.38e-11
+ mcm5m3l1_ca_w_2_400_s_2_100 = 4.70e-05  mcm5m3l1_cc_w_2_400_s_2_100 = 1.71e-11  mcm5m3l1_cf_w_2_400_s_2_100 = 3.59e-11
+ mcm5m3l1_ca_w_2_400_s_3_300 = 4.70e-05  mcm5m3l1_cc_w_2_400_s_3_300 = 6.29e-12  mcm5m3l1_cf_w_2_400_s_3_300 = 4.46e-11
+ mcm5m3l1_ca_w_2_400_s_9_000 = 4.70e-05  mcm5m3l1_cc_w_2_400_s_9_000 = 1.00e-13  mcm5m3l1_cf_w_2_400_s_9_000 = 5.04e-11
+ mcm5m3m1_ca_w_0_300_s_0_300 = 6.38e-05  mcm5m3m1_cc_w_0_300_s_0_300 = 1.07e-10  mcm5m3m1_cf_w_0_300_s_0_300 = 8.12e-12
+ mcm5m3m1_ca_w_0_300_s_0_360 = 6.38e-05  mcm5m3m1_cc_w_0_300_s_0_360 = 9.74e-11  mcm5m3m1_cf_w_0_300_s_0_360 = 9.86e-12
+ mcm5m3m1_ca_w_0_300_s_0_450 = 6.38e-05  mcm5m3m1_cc_w_0_300_s_0_450 = 8.50e-11  mcm5m3m1_cf_w_0_300_s_0_450 = 1.24e-11
+ mcm5m3m1_ca_w_0_300_s_0_600 = 6.38e-05  mcm5m3m1_cc_w_0_300_s_0_600 = 6.83e-11  mcm5m3m1_cf_w_0_300_s_0_600 = 1.65e-11
+ mcm5m3m1_ca_w_0_300_s_0_800 = 6.38e-05  mcm5m3m1_cc_w_0_300_s_0_800 = 5.25e-11  mcm5m3m1_cf_w_0_300_s_0_800 = 2.15e-11
+ mcm5m3m1_ca_w_0_300_s_1_000 = 6.38e-05  mcm5m3m1_cc_w_0_300_s_1_000 = 4.07e-11  mcm5m3m1_cf_w_0_300_s_1_000 = 2.61e-11
+ mcm5m3m1_ca_w_0_300_s_1_200 = 6.38e-05  mcm5m3m1_cc_w_0_300_s_1_200 = 3.20e-11  mcm5m3m1_cf_w_0_300_s_1_200 = 3.02e-11
+ mcm5m3m1_ca_w_0_300_s_2_100 = 6.38e-05  mcm5m3m1_cc_w_0_300_s_2_100 = 1.23e-11  mcm5m3m1_cf_w_0_300_s_2_100 = 4.30e-11
+ mcm5m3m1_ca_w_0_300_s_3_300 = 6.38e-05  mcm5m3m1_cc_w_0_300_s_3_300 = 3.77e-12  mcm5m3m1_cf_w_0_300_s_3_300 = 5.03e-11
+ mcm5m3m1_ca_w_0_300_s_9_000 = 6.38e-05  mcm5m3m1_cc_w_0_300_s_9_000 = 3.50e-14  mcm5m3m1_cf_w_0_300_s_9_000 = 5.40e-11
+ mcm5m3m1_ca_w_2_400_s_0_300 = 6.38e-05  mcm5m3m1_cc_w_2_400_s_0_300 = 1.13e-10  mcm5m3m1_cf_w_2_400_s_0_300 = 8.13e-12
+ mcm5m3m1_ca_w_2_400_s_0_360 = 6.38e-05  mcm5m3m1_cc_w_2_400_s_0_360 = 1.02e-10  mcm5m3m1_cf_w_2_400_s_0_360 = 9.88e-12
+ mcm5m3m1_ca_w_2_400_s_0_450 = 6.38e-05  mcm5m3m1_cc_w_2_400_s_0_450 = 8.90e-11  mcm5m3m1_cf_w_2_400_s_0_450 = 1.24e-11
+ mcm5m3m1_ca_w_2_400_s_0_600 = 6.38e-05  mcm5m3m1_cc_w_2_400_s_0_600 = 7.16e-11  mcm5m3m1_cf_w_2_400_s_0_600 = 1.65e-11
+ mcm5m3m1_ca_w_2_400_s_0_800 = 6.38e-05  mcm5m3m1_cc_w_2_400_s_0_800 = 5.50e-11  mcm5m3m1_cf_w_2_400_s_0_800 = 2.16e-11
+ mcm5m3m1_ca_w_2_400_s_1_000 = 6.38e-05  mcm5m3m1_cc_w_2_400_s_1_000 = 4.27e-11  mcm5m3m1_cf_w_2_400_s_1_000 = 2.63e-11
+ mcm5m3m1_ca_w_2_400_s_1_200 = 6.38e-05  mcm5m3m1_cc_w_2_400_s_1_200 = 3.36e-11  mcm5m3m1_cf_w_2_400_s_1_200 = 3.04e-11
+ mcm5m3m1_ca_w_2_400_s_2_100 = 6.38e-05  mcm5m3m1_cc_w_2_400_s_2_100 = 1.30e-11  mcm5m3m1_cf_w_2_400_s_2_100 = 4.35e-11
+ mcm5m3m1_ca_w_2_400_s_3_300 = 6.38e-05  mcm5m3m1_cc_w_2_400_s_3_300 = 4.01e-12  mcm5m3m1_cf_w_2_400_s_3_300 = 5.13e-11
+ mcm5m3m1_ca_w_2_400_s_9_000 = 6.38e-05  mcm5m3m1_cc_w_2_400_s_9_000 = 5.00e-14  mcm5m3m1_cf_w_2_400_s_9_000 = 5.51e-11
+ mcm5m3m2_ca_w_0_300_s_0_300 = 1.35e-04  mcm5m3m2_cc_w_0_300_s_0_300 = 9.76e-11  mcm5m3m2_cf_w_0_300_s_0_300 = 1.61e-11
+ mcm5m3m2_ca_w_0_300_s_0_360 = 1.35e-04  mcm5m3m2_cc_w_0_300_s_0_360 = 8.76e-11  mcm5m3m2_cf_w_0_300_s_0_360 = 1.93e-11
+ mcm5m3m2_ca_w_0_300_s_0_450 = 1.35e-04  mcm5m3m2_cc_w_0_300_s_0_450 = 7.54e-11  mcm5m3m2_cf_w_0_300_s_0_450 = 2.37e-11
+ mcm5m3m2_ca_w_0_300_s_0_600 = 1.35e-04  mcm5m3m2_cc_w_0_300_s_0_600 = 5.89e-11  mcm5m3m2_cf_w_0_300_s_0_600 = 3.02e-11
+ mcm5m3m2_ca_w_0_300_s_0_800 = 1.35e-04  mcm5m3m2_cc_w_0_300_s_0_800 = 4.35e-11  mcm5m3m2_cf_w_0_300_s_0_800 = 3.75e-11
+ mcm5m3m2_ca_w_0_300_s_1_000 = 1.35e-04  mcm5m3m2_cc_w_0_300_s_1_000 = 3.22e-11  mcm5m3m2_cf_w_0_300_s_1_000 = 4.36e-11
+ mcm5m3m2_ca_w_0_300_s_1_200 = 1.35e-04  mcm5m3m2_cc_w_0_300_s_1_200 = 2.43e-11  mcm5m3m2_cf_w_0_300_s_1_200 = 4.84e-11
+ mcm5m3m2_ca_w_0_300_s_2_100 = 1.35e-04  mcm5m3m2_cc_w_0_300_s_2_100 = 7.74e-12  mcm5m3m2_cf_w_0_300_s_2_100 = 6.13e-11
+ mcm5m3m2_ca_w_0_300_s_3_300 = 1.35e-04  mcm5m3m2_cc_w_0_300_s_3_300 = 1.85e-12  mcm5m3m2_cf_w_0_300_s_3_300 = 6.67e-11
+ mcm5m3m2_ca_w_0_300_s_9_000 = 1.35e-04  mcm5m3m2_cc_w_0_300_s_9_000 = 7.00e-14  mcm5m3m2_cf_w_0_300_s_9_000 = 6.88e-11
+ mcm5m3m2_ca_w_2_400_s_0_300 = 1.35e-04  mcm5m3m2_cc_w_2_400_s_0_300 = 1.02e-10  mcm5m3m2_cf_w_2_400_s_0_300 = 1.61e-11
+ mcm5m3m2_ca_w_2_400_s_0_360 = 1.35e-04  mcm5m3m2_cc_w_2_400_s_0_360 = 9.16e-11  mcm5m3m2_cf_w_2_400_s_0_360 = 1.93e-11
+ mcm5m3m2_ca_w_2_400_s_0_450 = 1.35e-04  mcm5m3m2_cc_w_2_400_s_0_450 = 7.84e-11  mcm5m3m2_cf_w_2_400_s_0_450 = 2.37e-11
+ mcm5m3m2_ca_w_2_400_s_0_600 = 1.35e-04  mcm5m3m2_cc_w_2_400_s_0_600 = 6.15e-11  mcm5m3m2_cf_w_2_400_s_0_600 = 3.02e-11
+ mcm5m3m2_ca_w_2_400_s_0_800 = 1.35e-04  mcm5m3m2_cc_w_2_400_s_0_800 = 4.55e-11  mcm5m3m2_cf_w_2_400_s_0_800 = 3.76e-11
+ mcm5m3m2_ca_w_2_400_s_1_000 = 1.35e-04  mcm5m3m2_cc_w_2_400_s_1_000 = 3.40e-11  mcm5m3m2_cf_w_2_400_s_1_000 = 4.37e-11
+ mcm5m3m2_ca_w_2_400_s_1_200 = 1.35e-04  mcm5m3m2_cc_w_2_400_s_1_200 = 2.56e-11  mcm5m3m2_cf_w_2_400_s_1_200 = 4.86e-11
+ mcm5m3m2_ca_w_2_400_s_2_100 = 1.35e-04  mcm5m3m2_cc_w_2_400_s_2_100 = 8.26e-12  mcm5m3m2_cf_w_2_400_s_2_100 = 6.18e-11
+ mcm5m3m2_ca_w_2_400_s_3_300 = 1.35e-04  mcm5m3m2_cc_w_2_400_s_3_300 = 2.07e-12  mcm5m3m2_cf_w_2_400_s_3_300 = 6.77e-11
+ mcm5m3m2_ca_w_2_400_s_9_000 = 1.35e-04  mcm5m3m2_cc_w_2_400_s_9_000 = 7.00e-14  mcm5m3m2_cf_w_2_400_s_9_000 = 6.98e-11
+ mcrdlm3f_ca_w_0_300_s_0_300 = 1.96e-05  mcrdlm3f_cc_w_0_300_s_0_300 = 1.17e-10  mcrdlm3f_cf_w_0_300_s_0_300 = 2.58e-12
+ mcrdlm3f_ca_w_0_300_s_0_360 = 1.96e-05  mcrdlm3f_cc_w_0_300_s_0_360 = 1.08e-10  mcrdlm3f_cf_w_0_300_s_0_360 = 3.16e-12
+ mcrdlm3f_ca_w_0_300_s_0_450 = 1.96e-05  mcrdlm3f_cc_w_0_300_s_0_450 = 9.65e-11  mcrdlm3f_cf_w_0_300_s_0_450 = 4.03e-12
+ mcrdlm3f_ca_w_0_300_s_0_600 = 1.96e-05  mcrdlm3f_cc_w_0_300_s_0_600 = 8.19e-11  mcrdlm3f_cf_w_0_300_s_0_600 = 5.47e-12
+ mcrdlm3f_ca_w_0_300_s_0_800 = 1.96e-05  mcrdlm3f_cc_w_0_300_s_0_800 = 6.73e-11  mcrdlm3f_cf_w_0_300_s_0_800 = 7.19e-12
+ mcrdlm3f_ca_w_0_300_s_1_000 = 1.96e-05  mcrdlm3f_cc_w_0_300_s_1_000 = 5.68e-11  mcrdlm3f_cf_w_0_300_s_1_000 = 8.95e-12
+ mcrdlm3f_ca_w_0_300_s_1_200 = 1.96e-05  mcrdlm3f_cc_w_0_300_s_1_200 = 4.89e-11  mcrdlm3f_cf_w_0_300_s_1_200 = 1.06e-11
+ mcrdlm3f_ca_w_0_300_s_2_100 = 1.96e-05  mcrdlm3f_cc_w_0_300_s_2_100 = 2.93e-11  mcrdlm3f_cf_w_0_300_s_2_100 = 1.76e-11
+ mcrdlm3f_ca_w_0_300_s_3_300 = 1.96e-05  mcrdlm3f_cc_w_0_300_s_3_300 = 1.76e-11  mcrdlm3f_cf_w_0_300_s_3_300 = 2.41e-11
+ mcrdlm3f_ca_w_0_300_s_9_000 = 1.96e-05  mcrdlm3f_cc_w_0_300_s_9_000 = 2.53e-12  mcrdlm3f_cf_w_0_300_s_9_000 = 3.62e-11
+ mcrdlm3f_ca_w_2_400_s_0_300 = 1.96e-05  mcrdlm3f_cc_w_2_400_s_0_300 = 1.37e-10  mcrdlm3f_cf_w_2_400_s_0_300 = 2.64e-12
+ mcrdlm3f_ca_w_2_400_s_0_360 = 1.96e-05  mcrdlm3f_cc_w_2_400_s_0_360 = 1.27e-10  mcrdlm3f_cf_w_2_400_s_0_360 = 3.21e-12
+ mcrdlm3f_ca_w_2_400_s_0_450 = 1.96e-05  mcrdlm3f_cc_w_2_400_s_0_450 = 1.14e-10  mcrdlm3f_cf_w_2_400_s_0_450 = 4.06e-12
+ mcrdlm3f_ca_w_2_400_s_0_600 = 1.96e-05  mcrdlm3f_cc_w_2_400_s_0_600 = 9.69e-11  mcrdlm3f_cf_w_2_400_s_0_600 = 5.45e-12
+ mcrdlm3f_ca_w_2_400_s_0_800 = 1.96e-05  mcrdlm3f_cc_w_2_400_s_0_800 = 8.03e-11  mcrdlm3f_cf_w_2_400_s_0_800 = 7.27e-12
+ mcrdlm3f_ca_w_2_400_s_1_000 = 1.96e-05  mcrdlm3f_cc_w_2_400_s_1_000 = 6.81e-11  mcrdlm3f_cf_w_2_400_s_1_000 = 9.05e-12
+ mcrdlm3f_ca_w_2_400_s_1_200 = 1.96e-05  mcrdlm3f_cc_w_2_400_s_1_200 = 5.89e-11  mcrdlm3f_cf_w_2_400_s_1_200 = 1.08e-11
+ mcrdlm3f_ca_w_2_400_s_2_100 = 1.96e-05  mcrdlm3f_cc_w_2_400_s_2_100 = 3.61e-11  mcrdlm3f_cf_w_2_400_s_2_100 = 1.77e-11
+ mcrdlm3f_ca_w_2_400_s_3_300 = 1.96e-05  mcrdlm3f_cc_w_2_400_s_3_300 = 2.21e-11  mcrdlm3f_cf_w_2_400_s_3_300 = 2.49e-11
+ mcrdlm3f_ca_w_2_400_s_9_000 = 1.96e-05  mcrdlm3f_cc_w_2_400_s_9_000 = 3.41e-12  mcrdlm3f_cf_w_2_400_s_9_000 = 3.93e-11
+ mcrdlm3d_ca_w_0_300_s_0_300 = 2.13e-05  mcrdlm3d_cc_w_0_300_s_0_300 = 1.17e-10  mcrdlm3d_cf_w_0_300_s_0_300 = 2.81e-12
+ mcrdlm3d_ca_w_0_300_s_0_360 = 2.13e-05  mcrdlm3d_cc_w_0_300_s_0_360 = 1.08e-10  mcrdlm3d_cf_w_0_300_s_0_360 = 3.43e-12
+ mcrdlm3d_ca_w_0_300_s_0_450 = 2.13e-05  mcrdlm3d_cc_w_0_300_s_0_450 = 9.60e-11  mcrdlm3d_cf_w_0_300_s_0_450 = 4.37e-12
+ mcrdlm3d_ca_w_0_300_s_0_600 = 2.13e-05  mcrdlm3d_cc_w_0_300_s_0_600 = 8.14e-11  mcrdlm3d_cf_w_0_300_s_0_600 = 5.92e-12
+ mcrdlm3d_ca_w_0_300_s_0_800 = 2.13e-05  mcrdlm3d_cc_w_0_300_s_0_800 = 6.67e-11  mcrdlm3d_cf_w_0_300_s_0_800 = 7.78e-12
+ mcrdlm3d_ca_w_0_300_s_1_000 = 2.13e-05  mcrdlm3d_cc_w_0_300_s_1_000 = 5.61e-11  mcrdlm3d_cf_w_0_300_s_1_000 = 9.68e-12
+ mcrdlm3d_ca_w_0_300_s_1_200 = 2.13e-05  mcrdlm3d_cc_w_0_300_s_1_200 = 4.82e-11  mcrdlm3d_cf_w_0_300_s_1_200 = 1.15e-11
+ mcrdlm3d_ca_w_0_300_s_2_100 = 2.13e-05  mcrdlm3d_cc_w_0_300_s_2_100 = 2.83e-11  mcrdlm3d_cf_w_0_300_s_2_100 = 1.88e-11
+ mcrdlm3d_ca_w_0_300_s_3_300 = 2.13e-05  mcrdlm3d_cc_w_0_300_s_3_300 = 1.67e-11  mcrdlm3d_cf_w_0_300_s_3_300 = 2.55e-11
+ mcrdlm3d_ca_w_0_300_s_9_000 = 2.13e-05  mcrdlm3d_cc_w_0_300_s_9_000 = 2.27e-12  mcrdlm3d_cf_w_0_300_s_9_000 = 3.74e-11
+ mcrdlm3d_ca_w_2_400_s_0_300 = 2.13e-05  mcrdlm3d_cc_w_2_400_s_0_300 = 1.36e-10  mcrdlm3d_cf_w_2_400_s_0_300 = 2.87e-12
+ mcrdlm3d_ca_w_2_400_s_0_360 = 2.13e-05  mcrdlm3d_cc_w_2_400_s_0_360 = 1.26e-10  mcrdlm3d_cf_w_2_400_s_0_360 = 3.49e-12
+ mcrdlm3d_ca_w_2_400_s_0_450 = 2.13e-05  mcrdlm3d_cc_w_2_400_s_0_450 = 1.13e-10  mcrdlm3d_cf_w_2_400_s_0_450 = 4.41e-12
+ mcrdlm3d_ca_w_2_400_s_0_600 = 2.13e-05  mcrdlm3d_cc_w_2_400_s_0_600 = 9.58e-11  mcrdlm3d_cf_w_2_400_s_0_600 = 5.92e-12
+ mcrdlm3d_ca_w_2_400_s_0_800 = 2.13e-05  mcrdlm3d_cc_w_2_400_s_0_800 = 7.92e-11  mcrdlm3d_cf_w_2_400_s_0_800 = 7.88e-12
+ mcrdlm3d_ca_w_2_400_s_1_000 = 2.13e-05  mcrdlm3d_cc_w_2_400_s_1_000 = 6.70e-11  mcrdlm3d_cf_w_2_400_s_1_000 = 9.79e-12
+ mcrdlm3d_ca_w_2_400_s_1_200 = 2.13e-05  mcrdlm3d_cc_w_2_400_s_1_200 = 5.77e-11  mcrdlm3d_cf_w_2_400_s_1_200 = 1.16e-11
+ mcrdlm3d_ca_w_2_400_s_2_100 = 2.13e-05  mcrdlm3d_cc_w_2_400_s_2_100 = 3.50e-11  mcrdlm3d_cf_w_2_400_s_2_100 = 1.89e-11
+ mcrdlm3d_ca_w_2_400_s_3_300 = 2.13e-05  mcrdlm3d_cc_w_2_400_s_3_300 = 2.11e-11  mcrdlm3d_cf_w_2_400_s_3_300 = 2.64e-11
+ mcrdlm3d_ca_w_2_400_s_9_000 = 2.13e-05  mcrdlm3d_cc_w_2_400_s_9_000 = 3.11e-12  mcrdlm3d_cf_w_2_400_s_9_000 = 4.06e-11
+ mcrdlm3p1_ca_w_0_300_s_0_300 = 2.39e-05  mcrdlm3p1_cc_w_0_300_s_0_300 = 1.16e-10  mcrdlm3p1_cf_w_0_300_s_0_300 = 3.15e-12
+ mcrdlm3p1_ca_w_0_300_s_0_360 = 2.39e-05  mcrdlm3p1_cc_w_0_300_s_0_360 = 1.07e-10  mcrdlm3p1_cf_w_0_300_s_0_360 = 3.84e-12
+ mcrdlm3p1_ca_w_0_300_s_0_450 = 2.39e-05  mcrdlm3p1_cc_w_0_300_s_0_450 = 9.53e-11  mcrdlm3p1_cf_w_0_300_s_0_450 = 4.89e-12
+ mcrdlm3p1_ca_w_0_300_s_0_600 = 2.39e-05  mcrdlm3p1_cc_w_0_300_s_0_600 = 8.03e-11  mcrdlm3p1_cf_w_0_300_s_0_600 = 6.60e-12
+ mcrdlm3p1_ca_w_0_300_s_0_800 = 2.39e-05  mcrdlm3p1_cc_w_0_300_s_0_800 = 6.57e-11  mcrdlm3p1_cf_w_0_300_s_0_800 = 8.67e-12
+ mcrdlm3p1_ca_w_0_300_s_1_000 = 2.39e-05  mcrdlm3p1_cc_w_0_300_s_1_000 = 5.51e-11  mcrdlm3p1_cf_w_0_300_s_1_000 = 1.08e-11
+ mcrdlm3p1_ca_w_0_300_s_1_200 = 2.39e-05  mcrdlm3p1_cc_w_0_300_s_1_200 = 4.70e-11  mcrdlm3p1_cf_w_0_300_s_1_200 = 1.27e-11
+ mcrdlm3p1_ca_w_0_300_s_2_100 = 2.39e-05  mcrdlm3p1_cc_w_0_300_s_2_100 = 2.72e-11  mcrdlm3p1_cf_w_0_300_s_2_100 = 2.06e-11
+ mcrdlm3p1_ca_w_0_300_s_3_300 = 2.39e-05  mcrdlm3p1_cc_w_0_300_s_3_300 = 1.56e-11  mcrdlm3p1_cf_w_0_300_s_3_300 = 2.76e-11
+ mcrdlm3p1_ca_w_0_300_s_9_000 = 2.39e-05  mcrdlm3p1_cc_w_0_300_s_9_000 = 1.96e-12  mcrdlm3p1_cf_w_0_300_s_9_000 = 3.90e-11
+ mcrdlm3p1_ca_w_2_400_s_0_300 = 2.39e-05  mcrdlm3p1_cc_w_2_400_s_0_300 = 1.35e-10  mcrdlm3p1_cf_w_2_400_s_0_300 = 3.25e-12
+ mcrdlm3p1_ca_w_2_400_s_0_360 = 2.39e-05  mcrdlm3p1_cc_w_2_400_s_0_360 = 1.25e-10  mcrdlm3p1_cf_w_2_400_s_0_360 = 3.94e-12
+ mcrdlm3p1_ca_w_2_400_s_0_450 = 2.39e-05  mcrdlm3p1_cc_w_2_400_s_0_450 = 1.11e-10  mcrdlm3p1_cf_w_2_400_s_0_450 = 4.97e-12
+ mcrdlm3p1_ca_w_2_400_s_0_600 = 2.39e-05  mcrdlm3p1_cc_w_2_400_s_0_600 = 9.40e-11  mcrdlm3p1_cf_w_2_400_s_0_600 = 6.64e-12
+ mcrdlm3p1_ca_w_2_400_s_0_800 = 2.39e-05  mcrdlm3p1_cc_w_2_400_s_0_800 = 7.76e-11  mcrdlm3p1_cf_w_2_400_s_0_800 = 8.81e-12
+ mcrdlm3p1_ca_w_2_400_s_1_000 = 2.39e-05  mcrdlm3p1_cc_w_2_400_s_1_000 = 6.54e-11  mcrdlm3p1_cf_w_2_400_s_1_000 = 1.09e-11
+ mcrdlm3p1_ca_w_2_400_s_1_200 = 2.39e-05  mcrdlm3p1_cc_w_2_400_s_1_200 = 5.62e-11  mcrdlm3p1_cf_w_2_400_s_1_200 = 1.29e-11
+ mcrdlm3p1_ca_w_2_400_s_2_100 = 2.39e-05  mcrdlm3p1_cc_w_2_400_s_2_100 = 3.35e-11  mcrdlm3p1_cf_w_2_400_s_2_100 = 2.08e-11
+ mcrdlm3p1_ca_w_2_400_s_3_300 = 2.39e-05  mcrdlm3p1_cc_w_2_400_s_3_300 = 1.98e-11  mcrdlm3p1_cf_w_2_400_s_3_300 = 2.86e-11
+ mcrdlm3p1_ca_w_2_400_s_9_000 = 2.39e-05  mcrdlm3p1_cc_w_2_400_s_9_000 = 2.75e-12  mcrdlm3p1_cf_w_2_400_s_9_000 = 4.25e-11
+ mcrdlm3l1_ca_w_0_300_s_0_300 = 2.87e-05  mcrdlm3l1_cc_w_0_300_s_0_300 = 1.15e-10  mcrdlm3l1_cf_w_0_300_s_0_300 = 3.74e-12
+ mcrdlm3l1_ca_w_0_300_s_0_360 = 2.87e-05  mcrdlm3l1_cc_w_0_300_s_0_360 = 1.06e-10  mcrdlm3l1_cf_w_0_300_s_0_360 = 4.55e-12
+ mcrdlm3l1_ca_w_0_300_s_0_450 = 2.87e-05  mcrdlm3l1_cc_w_0_300_s_0_450 = 9.40e-11  mcrdlm3l1_cf_w_0_300_s_0_450 = 5.79e-12
+ mcrdlm3l1_ca_w_0_300_s_0_600 = 2.87e-05  mcrdlm3l1_cc_w_0_300_s_0_600 = 7.89e-11  mcrdlm3l1_cf_w_0_300_s_0_600 = 7.78e-12
+ mcrdlm3l1_ca_w_0_300_s_0_800 = 2.87e-05  mcrdlm3l1_cc_w_0_300_s_0_800 = 6.42e-11  mcrdlm3l1_cf_w_0_300_s_0_800 = 1.02e-11
+ mcrdlm3l1_ca_w_0_300_s_1_000 = 2.87e-05  mcrdlm3l1_cc_w_0_300_s_1_000 = 5.34e-11  mcrdlm3l1_cf_w_0_300_s_1_000 = 1.26e-11
+ mcrdlm3l1_ca_w_0_300_s_1_200 = 2.87e-05  mcrdlm3l1_cc_w_0_300_s_1_200 = 4.52e-11  mcrdlm3l1_cf_w_0_300_s_1_200 = 1.48e-11
+ mcrdlm3l1_ca_w_0_300_s_2_100 = 2.87e-05  mcrdlm3l1_cc_w_0_300_s_2_100 = 2.53e-11  mcrdlm3l1_cf_w_0_300_s_2_100 = 2.36e-11
+ mcrdlm3l1_ca_w_0_300_s_3_300 = 2.87e-05  mcrdlm3l1_cc_w_0_300_s_3_300 = 1.41e-11  mcrdlm3l1_cf_w_0_300_s_3_300 = 3.09e-11
+ mcrdlm3l1_ca_w_0_300_s_9_000 = 2.87e-05  mcrdlm3l1_cc_w_0_300_s_9_000 = 1.61e-12  mcrdlm3l1_cf_w_0_300_s_9_000 = 4.17e-11
+ mcrdlm3l1_ca_w_2_400_s_0_300 = 2.87e-05  mcrdlm3l1_cc_w_2_400_s_0_300 = 1.33e-10  mcrdlm3l1_cf_w_2_400_s_0_300 = 3.79e-12
+ mcrdlm3l1_ca_w_2_400_s_0_360 = 2.87e-05  mcrdlm3l1_cc_w_2_400_s_0_360 = 1.22e-10  mcrdlm3l1_cf_w_2_400_s_0_360 = 4.60e-12
+ mcrdlm3l1_ca_w_2_400_s_0_450 = 2.87e-05  mcrdlm3l1_cc_w_2_400_s_0_450 = 1.09e-10  mcrdlm3l1_cf_w_2_400_s_0_450 = 5.81e-12
+ mcrdlm3l1_ca_w_2_400_s_0_600 = 2.87e-05  mcrdlm3l1_cc_w_2_400_s_0_600 = 9.15e-11  mcrdlm3l1_cf_w_2_400_s_0_600 = 7.77e-12
+ mcrdlm3l1_ca_w_2_400_s_0_800 = 2.87e-05  mcrdlm3l1_cc_w_2_400_s_0_800 = 7.53e-11  mcrdlm3l1_cf_w_2_400_s_0_800 = 1.03e-11
+ mcrdlm3l1_ca_w_2_400_s_1_000 = 2.87e-05  mcrdlm3l1_cc_w_2_400_s_1_000 = 6.30e-11  mcrdlm3l1_cf_w_2_400_s_1_000 = 1.27e-11
+ mcrdlm3l1_ca_w_2_400_s_1_200 = 2.87e-05  mcrdlm3l1_cc_w_2_400_s_1_200 = 5.38e-11  mcrdlm3l1_cf_w_2_400_s_1_200 = 1.50e-11
+ mcrdlm3l1_ca_w_2_400_s_2_100 = 2.87e-05  mcrdlm3l1_cc_w_2_400_s_2_100 = 3.15e-11  mcrdlm3l1_cf_w_2_400_s_2_100 = 2.37e-11
+ mcrdlm3l1_ca_w_2_400_s_3_300 = 2.87e-05  mcrdlm3l1_cc_w_2_400_s_3_300 = 1.81e-11  mcrdlm3l1_cf_w_2_400_s_3_300 = 3.19e-11
+ mcrdlm3l1_ca_w_2_400_s_9_000 = 2.87e-05  mcrdlm3l1_cc_w_2_400_s_9_000 = 2.30e-12  mcrdlm3l1_cf_w_2_400_s_9_000 = 4.51e-11
+ mcrdlm3m1_ca_w_0_300_s_0_300 = 4.55e-05  mcrdlm3m1_cc_w_0_300_s_0_300 = 1.12e-10  mcrdlm3m1_cf_w_0_300_s_0_300 = 5.82e-12
+ mcrdlm3m1_ca_w_0_300_s_0_360 = 4.55e-05  mcrdlm3m1_cc_w_0_300_s_0_360 = 1.02e-10  mcrdlm3m1_cf_w_0_300_s_0_360 = 7.05e-12
+ mcrdlm3m1_ca_w_0_300_s_0_450 = 4.55e-05  mcrdlm3m1_cc_w_0_300_s_0_450 = 9.01e-11  mcrdlm3m1_cf_w_0_300_s_0_450 = 8.88e-12
+ mcrdlm3m1_ca_w_0_300_s_0_600 = 4.55e-05  mcrdlm3m1_cc_w_0_300_s_0_600 = 7.44e-11  mcrdlm3m1_cf_w_0_300_s_0_600 = 1.18e-11
+ mcrdlm3m1_ca_w_0_300_s_0_800 = 4.55e-05  mcrdlm3m1_cc_w_0_300_s_0_800 = 5.96e-11  mcrdlm3m1_cf_w_0_300_s_0_800 = 1.53e-11
+ mcrdlm3m1_ca_w_0_300_s_1_000 = 4.55e-05  mcrdlm3m1_cc_w_0_300_s_1_000 = 4.87e-11  mcrdlm3m1_cf_w_0_300_s_1_000 = 1.86e-11
+ mcrdlm3m1_ca_w_0_300_s_1_200 = 4.55e-05  mcrdlm3m1_cc_w_0_300_s_1_200 = 4.07e-11  mcrdlm3m1_cf_w_0_300_s_1_200 = 2.16e-11
+ mcrdlm3m1_ca_w_0_300_s_2_100 = 4.55e-05  mcrdlm3m1_cc_w_0_300_s_2_100 = 2.09e-11  mcrdlm3m1_cf_w_0_300_s_2_100 = 3.22e-11
+ mcrdlm3m1_ca_w_0_300_s_3_300 = 4.55e-05  mcrdlm3m1_cc_w_0_300_s_3_300 = 1.08e-11  mcrdlm3m1_cf_w_0_300_s_3_300 = 3.99e-11
+ mcrdlm3m1_ca_w_0_300_s_9_000 = 4.55e-05  mcrdlm3m1_cc_w_0_300_s_9_000 = 1.06e-12  mcrdlm3m1_cf_w_0_300_s_9_000 = 4.87e-11
+ mcrdlm3m1_ca_w_2_400_s_0_300 = 4.55e-05  mcrdlm3m1_cc_w_2_400_s_0_300 = 1.27e-10  mcrdlm3m1_cf_w_2_400_s_0_300 = 5.82e-12
+ mcrdlm3m1_ca_w_2_400_s_0_360 = 4.55e-05  mcrdlm3m1_cc_w_2_400_s_0_360 = 1.17e-10  mcrdlm3m1_cf_w_2_400_s_0_360 = 7.06e-12
+ mcrdlm3m1_ca_w_2_400_s_0_450 = 4.55e-05  mcrdlm3m1_cc_w_2_400_s_0_450 = 1.03e-10  mcrdlm3m1_cf_w_2_400_s_0_450 = 8.88e-12
+ mcrdlm3m1_ca_w_2_400_s_0_600 = 4.55e-05  mcrdlm3m1_cc_w_2_400_s_0_600 = 8.58e-11  mcrdlm3m1_cf_w_2_400_s_0_600 = 1.18e-11
+ mcrdlm3m1_ca_w_2_400_s_0_800 = 4.55e-05  mcrdlm3m1_cc_w_2_400_s_0_800 = 6.96e-11  mcrdlm3m1_cf_w_2_400_s_0_800 = 1.54e-11
+ mcrdlm3m1_ca_w_2_400_s_1_000 = 4.55e-05  mcrdlm3m1_cc_w_2_400_s_1_000 = 5.75e-11  mcrdlm3m1_cf_w_2_400_s_1_000 = 1.87e-11
+ mcrdlm3m1_ca_w_2_400_s_1_200 = 4.55e-05  mcrdlm3m1_cc_w_2_400_s_1_200 = 4.85e-11  mcrdlm3m1_cf_w_2_400_s_1_200 = 2.17e-11
+ mcrdlm3m1_ca_w_2_400_s_2_100 = 4.55e-05  mcrdlm3m1_cc_w_2_400_s_2_100 = 2.68e-11  mcrdlm3m1_cf_w_2_400_s_2_100 = 3.23e-11
+ mcrdlm3m1_ca_w_2_400_s_3_300 = 4.55e-05  mcrdlm3m1_cc_w_2_400_s_3_300 = 1.46e-11  mcrdlm3m1_cf_w_2_400_s_3_300 = 4.10e-11
+ mcrdlm3m1_ca_w_2_400_s_9_000 = 4.55e-05  mcrdlm3m1_cc_w_2_400_s_9_000 = 1.60e-12  mcrdlm3m1_cf_w_2_400_s_9_000 = 5.26e-11
+ mcrdlm3m2_ca_w_0_300_s_0_300 = 1.17e-04  mcrdlm3m2_cc_w_0_300_s_0_300 = 1.02e-10  mcrdlm3m2_cf_w_0_300_s_0_300 = 1.38e-11
+ mcrdlm3m2_ca_w_0_300_s_0_360 = 1.17e-04  mcrdlm3m2_cc_w_0_300_s_0_360 = 9.27e-11  mcrdlm3m2_cf_w_0_300_s_0_360 = 1.65e-11
+ mcrdlm3m2_ca_w_0_300_s_0_450 = 1.17e-04  mcrdlm3m2_cc_w_0_300_s_0_450 = 8.04e-11  mcrdlm3m2_cf_w_0_300_s_0_450 = 2.01e-11
+ mcrdlm3m2_ca_w_0_300_s_0_600 = 1.17e-04  mcrdlm3m2_cc_w_0_300_s_0_600 = 6.51e-11  mcrdlm3m2_cf_w_0_300_s_0_600 = 2.55e-11
+ mcrdlm3m2_ca_w_0_300_s_0_800 = 1.17e-04  mcrdlm3m2_cc_w_0_300_s_0_800 = 5.07e-11  mcrdlm3m2_cf_w_0_300_s_0_800 = 3.14e-11
+ mcrdlm3m2_ca_w_0_300_s_1_000 = 1.17e-04  mcrdlm3m2_cc_w_0_300_s_1_000 = 4.01e-11  mcrdlm3m2_cf_w_0_300_s_1_000 = 3.63e-11
+ mcrdlm3m2_ca_w_0_300_s_1_200 = 1.17e-04  mcrdlm3m2_cc_w_0_300_s_1_200 = 3.25e-11  mcrdlm3m2_cf_w_0_300_s_1_200 = 4.04e-11
+ mcrdlm3m2_ca_w_0_300_s_2_100 = 1.17e-04  mcrdlm3m2_cc_w_0_300_s_2_100 = 1.50e-11  mcrdlm3m2_cf_w_0_300_s_2_100 = 5.25e-11
+ mcrdlm3m2_ca_w_0_300_s_3_300 = 1.17e-04  mcrdlm3m2_cc_w_0_300_s_3_300 = 7.08e-12  mcrdlm3m2_cf_w_0_300_s_3_300 = 5.93e-11
+ mcrdlm3m2_ca_w_0_300_s_9_000 = 1.17e-04  mcrdlm3m2_cc_w_0_300_s_9_000 = 5.55e-13  mcrdlm3m2_cf_w_0_300_s_9_000 = 6.56e-11
+ mcrdlm3m2_ca_w_2_400_s_0_300 = 1.17e-04  mcrdlm3m2_cc_w_2_400_s_0_300 = 1.16e-10  mcrdlm3m2_cf_w_2_400_s_0_300 = 1.38e-11
+ mcrdlm3m2_ca_w_2_400_s_0_360 = 1.17e-04  mcrdlm3m2_cc_w_2_400_s_0_360 = 1.06e-10  mcrdlm3m2_cf_w_2_400_s_0_360 = 1.64e-11
+ mcrdlm3m2_ca_w_2_400_s_0_450 = 1.17e-04  mcrdlm3m2_cc_w_2_400_s_0_450 = 9.24e-11  mcrdlm3m2_cf_w_2_400_s_0_450 = 2.01e-11
+ mcrdlm3m2_ca_w_2_400_s_0_600 = 1.17e-04  mcrdlm3m2_cc_w_2_400_s_0_600 = 7.60e-11  mcrdlm3m2_cf_w_2_400_s_0_600 = 2.54e-11
+ mcrdlm3m2_ca_w_2_400_s_0_800 = 1.17e-04  mcrdlm3m2_cc_w_2_400_s_0_800 = 6.01e-11  mcrdlm3m2_cf_w_2_400_s_0_800 = 3.14e-11
+ mcrdlm3m2_ca_w_2_400_s_1_000 = 1.17e-04  mcrdlm3m2_cc_w_2_400_s_1_000 = 4.85e-11  mcrdlm3m2_cf_w_2_400_s_1_000 = 3.64e-11
+ mcrdlm3m2_ca_w_2_400_s_1_200 = 1.17e-04  mcrdlm3m2_cc_w_2_400_s_1_200 = 4.03e-11  mcrdlm3m2_cf_w_2_400_s_1_200 = 4.05e-11
+ mcrdlm3m2_ca_w_2_400_s_2_100 = 1.17e-04  mcrdlm3m2_cc_w_2_400_s_2_100 = 2.09e-11  mcrdlm3m2_cf_w_2_400_s_2_100 = 5.28e-11
+ mcrdlm3m2_ca_w_2_400_s_3_300 = 1.17e-04  mcrdlm3m2_cc_w_2_400_s_3_300 = 1.08e-11  mcrdlm3m2_cf_w_2_400_s_3_300 = 6.11e-11
+ mcrdlm3m2_ca_w_2_400_s_9_000 = 1.17e-04  mcrdlm3m2_cc_w_2_400_s_9_000 = 9.95e-13  mcrdlm3m2_cf_w_2_400_s_9_000 = 7.03e-11
+ mcm5m4f_ca_w_0_300_s_0_300 = 1.06e-04  mcm5m4f_cc_w_0_300_s_0_300 = 1.02e-10  mcm5m4f_cf_w_0_300_s_0_300 = 1.20e-11
+ mcm5m4f_ca_w_0_300_s_0_360 = 1.06e-04  mcm5m4f_cc_w_0_300_s_0_360 = 9.31e-11  mcm5m4f_cf_w_0_300_s_0_360 = 1.44e-11
+ mcm5m4f_ca_w_0_300_s_0_450 = 1.06e-04  mcm5m4f_cc_w_0_300_s_0_450 = 8.12e-11  mcm5m4f_cf_w_0_300_s_0_450 = 1.78e-11
+ mcm5m4f_ca_w_0_300_s_0_600 = 1.06e-04  mcm5m4f_cc_w_0_300_s_0_600 = 6.51e-11  mcm5m4f_cf_w_0_300_s_0_600 = 2.29e-11
+ mcm5m4f_ca_w_0_300_s_0_800 = 1.06e-04  mcm5m4f_cc_w_0_300_s_0_800 = 4.99e-11  mcm5m4f_cf_w_0_300_s_0_800 = 2.87e-11
+ mcm5m4f_ca_w_0_300_s_1_000 = 1.06e-04  mcm5m4f_cc_w_0_300_s_1_000 = 3.90e-11  mcm5m4f_cf_w_0_300_s_1_000 = 3.37e-11
+ mcm5m4f_ca_w_0_300_s_1_200 = 1.06e-04  mcm5m4f_cc_w_0_300_s_1_200 = 3.10e-11  mcm5m4f_cf_w_0_300_s_1_200 = 3.79e-11
+ mcm5m4f_ca_w_0_300_s_2_100 = 1.06e-04  mcm5m4f_cc_w_0_300_s_2_100 = 1.29e-11  mcm5m4f_cf_w_0_300_s_2_100 = 5.01e-11
+ mcm5m4f_ca_w_0_300_s_3_300 = 1.06e-04  mcm5m4f_cc_w_0_300_s_3_300 = 4.90e-12  mcm5m4f_cf_w_0_300_s_3_300 = 5.71e-11
+ mcm5m4f_ca_w_0_300_s_9_000 = 1.06e-04  mcm5m4f_cc_w_0_300_s_9_000 = 1.00e-13  mcm5m4f_cf_w_0_300_s_9_000 = 6.17e-11
+ mcm5m4f_ca_w_2_400_s_0_300 = 1.06e-04  mcm5m4f_cc_w_2_400_s_0_300 = 1.12e-10  mcm5m4f_cf_w_2_400_s_0_300 = 1.20e-11
+ mcm5m4f_ca_w_2_400_s_0_360 = 1.06e-04  mcm5m4f_cc_w_2_400_s_0_360 = 1.02e-10  mcm5m4f_cf_w_2_400_s_0_360 = 1.44e-11
+ mcm5m4f_ca_w_2_400_s_0_450 = 1.06e-04  mcm5m4f_cc_w_2_400_s_0_450 = 8.85e-11  mcm5m4f_cf_w_2_400_s_0_450 = 1.78e-11
+ mcm5m4f_ca_w_2_400_s_0_600 = 1.06e-04  mcm5m4f_cc_w_2_400_s_0_600 = 7.19e-11  mcm5m4f_cf_w_2_400_s_0_600 = 2.28e-11
+ mcm5m4f_ca_w_2_400_s_0_800 = 1.06e-04  mcm5m4f_cc_w_2_400_s_0_800 = 5.54e-11  mcm5m4f_cf_w_2_400_s_0_800 = 2.87e-11
+ mcm5m4f_ca_w_2_400_s_1_000 = 1.06e-04  mcm5m4f_cc_w_2_400_s_1_000 = 4.36e-11  mcm5m4f_cf_w_2_400_s_1_000 = 3.38e-11
+ mcm5m4f_ca_w_2_400_s_1_200 = 1.06e-04  mcm5m4f_cc_w_2_400_s_1_200 = 3.50e-11  mcm5m4f_cf_w_2_400_s_1_200 = 3.80e-11
+ mcm5m4f_ca_w_2_400_s_2_100 = 1.06e-04  mcm5m4f_cc_w_2_400_s_2_100 = 1.55e-11  mcm5m4f_cf_w_2_400_s_2_100 = 5.06e-11
+ mcm5m4f_ca_w_2_400_s_3_300 = 1.06e-04  mcm5m4f_cc_w_2_400_s_3_300 = 6.21e-12  mcm5m4f_cf_w_2_400_s_3_300 = 5.86e-11
+ mcm5m4f_ca_w_2_400_s_9_000 = 1.06e-04  mcm5m4f_cc_w_2_400_s_9_000 = 1.20e-13  mcm5m4f_cf_w_2_400_s_9_000 = 6.43e-11
+ mcm5m4d_ca_w_0_300_s_0_300 = 1.07e-04  mcm5m4d_cc_w_0_300_s_0_300 = 1.02e-10  mcm5m4d_cf_w_0_300_s_0_300 = 1.21e-11
+ mcm5m4d_ca_w_0_300_s_0_360 = 1.07e-04  mcm5m4d_cc_w_0_300_s_0_360 = 9.29e-11  mcm5m4d_cf_w_0_300_s_0_360 = 1.45e-11
+ mcm5m4d_ca_w_0_300_s_0_450 = 1.07e-04  mcm5m4d_cc_w_0_300_s_0_450 = 8.10e-11  mcm5m4d_cf_w_0_300_s_0_450 = 1.79e-11
+ mcm5m4d_ca_w_0_300_s_0_600 = 1.07e-04  mcm5m4d_cc_w_0_300_s_0_600 = 6.48e-11  mcm5m4d_cf_w_0_300_s_0_600 = 2.31e-11
+ mcm5m4d_ca_w_0_300_s_0_800 = 1.07e-04  mcm5m4d_cc_w_0_300_s_0_800 = 4.96e-11  mcm5m4d_cf_w_0_300_s_0_800 = 2.89e-11
+ mcm5m4d_ca_w_0_300_s_1_000 = 1.07e-04  mcm5m4d_cc_w_0_300_s_1_000 = 3.86e-11  mcm5m4d_cf_w_0_300_s_1_000 = 3.40e-11
+ mcm5m4d_ca_w_0_300_s_1_200 = 1.07e-04  mcm5m4d_cc_w_0_300_s_1_200 = 3.06e-11  mcm5m4d_cf_w_0_300_s_1_200 = 3.82e-11
+ mcm5m4d_ca_w_0_300_s_2_100 = 1.07e-04  mcm5m4d_cc_w_0_300_s_2_100 = 1.26e-11  mcm5m4d_cf_w_0_300_s_2_100 = 5.05e-11
+ mcm5m4d_ca_w_0_300_s_3_300 = 1.07e-04  mcm5m4d_cc_w_0_300_s_3_300 = 4.66e-12  mcm5m4d_cf_w_0_300_s_3_300 = 5.74e-11
+ mcm5m4d_ca_w_0_300_s_9_000 = 1.07e-04  mcm5m4d_cc_w_0_300_s_9_000 = 1.15e-13  mcm5m4d_cf_w_0_300_s_9_000 = 6.18e-11
+ mcm5m4d_ca_w_2_400_s_0_300 = 1.07e-04  mcm5m4d_cc_w_2_400_s_0_300 = 1.11e-10  mcm5m4d_cf_w_2_400_s_0_300 = 1.21e-11
+ mcm5m4d_ca_w_2_400_s_0_360 = 1.07e-04  mcm5m4d_cc_w_2_400_s_0_360 = 1.01e-10  mcm5m4d_cf_w_2_400_s_0_360 = 1.45e-11
+ mcm5m4d_ca_w_2_400_s_0_450 = 1.07e-04  mcm5m4d_cc_w_2_400_s_0_450 = 8.79e-11  mcm5m4d_cf_w_2_400_s_0_450 = 1.79e-11
+ mcm5m4d_ca_w_2_400_s_0_600 = 1.07e-04  mcm5m4d_cc_w_2_400_s_0_600 = 7.12e-11  mcm5m4d_cf_w_2_400_s_0_600 = 2.30e-11
+ mcm5m4d_ca_w_2_400_s_0_800 = 1.07e-04  mcm5m4d_cc_w_2_400_s_0_800 = 5.47e-11  mcm5m4d_cf_w_2_400_s_0_800 = 2.90e-11
+ mcm5m4d_ca_w_2_400_s_1_000 = 1.07e-04  mcm5m4d_cc_w_2_400_s_1_000 = 4.29e-11  mcm5m4d_cf_w_2_400_s_1_000 = 3.41e-11
+ mcm5m4d_ca_w_2_400_s_1_200 = 1.07e-04  mcm5m4d_cc_w_2_400_s_1_200 = 3.43e-11  mcm5m4d_cf_w_2_400_s_1_200 = 3.84e-11
+ mcm5m4d_ca_w_2_400_s_2_100 = 1.07e-04  mcm5m4d_cc_w_2_400_s_2_100 = 1.49e-11  mcm5m4d_cf_w_2_400_s_2_100 = 5.11e-11
+ mcm5m4d_ca_w_2_400_s_3_300 = 1.07e-04  mcm5m4d_cc_w_2_400_s_3_300 = 5.78e-12  mcm5m4d_cf_w_2_400_s_3_300 = 5.88e-11
+ mcm5m4d_ca_w_2_400_s_9_000 = 1.07e-04  mcm5m4d_cc_w_2_400_s_9_000 = 1.00e-13  mcm5m4d_cf_w_2_400_s_9_000 = 6.43e-11
+ mcm5m4p1_ca_w_0_300_s_0_300 = 1.08e-04  mcm5m4p1_cc_w_0_300_s_0_300 = 1.02e-10  mcm5m4p1_cf_w_0_300_s_0_300 = 1.22e-11
+ mcm5m4p1_ca_w_0_300_s_0_360 = 1.08e-04  mcm5m4p1_cc_w_0_300_s_0_360 = 9.26e-11  mcm5m4p1_cf_w_0_300_s_0_360 = 1.47e-11
+ mcm5m4p1_ca_w_0_300_s_0_450 = 1.08e-04  mcm5m4p1_cc_w_0_300_s_0_450 = 8.07e-11  mcm5m4p1_cf_w_0_300_s_0_450 = 1.81e-11
+ mcm5m4p1_ca_w_0_300_s_0_600 = 1.08e-04  mcm5m4p1_cc_w_0_300_s_0_600 = 6.44e-11  mcm5m4p1_cf_w_0_300_s_0_600 = 2.34e-11
+ mcm5m4p1_ca_w_0_300_s_0_800 = 1.08e-04  mcm5m4p1_cc_w_0_300_s_0_800 = 4.92e-11  mcm5m4p1_cf_w_0_300_s_0_800 = 2.93e-11
+ mcm5m4p1_ca_w_0_300_s_1_000 = 1.08e-04  mcm5m4p1_cc_w_0_300_s_1_000 = 3.82e-11  mcm5m4p1_cf_w_0_300_s_1_000 = 3.44e-11
+ mcm5m4p1_ca_w_0_300_s_1_200 = 1.08e-04  mcm5m4p1_cc_w_0_300_s_1_200 = 3.01e-11  mcm5m4p1_cf_w_0_300_s_1_200 = 3.87e-11
+ mcm5m4p1_ca_w_0_300_s_2_100 = 1.08e-04  mcm5m4p1_cc_w_0_300_s_2_100 = 1.21e-11  mcm5m4p1_cf_w_0_300_s_2_100 = 5.11e-11
+ mcm5m4p1_ca_w_0_300_s_3_300 = 1.08e-04  mcm5m4p1_cc_w_0_300_s_3_300 = 4.31e-12  mcm5m4p1_cf_w_0_300_s_3_300 = 5.78e-11
+ mcm5m4p1_ca_w_0_300_s_9_000 = 1.08e-04  mcm5m4p1_cc_w_0_300_s_9_000 = 6.50e-14  mcm5m4p1_cf_w_0_300_s_9_000 = 6.20e-11
+ mcm5m4p1_ca_w_2_400_s_0_300 = 1.08e-04  mcm5m4p1_cc_w_2_400_s_0_300 = 1.11e-10  mcm5m4p1_cf_w_2_400_s_0_300 = 1.23e-11
+ mcm5m4p1_ca_w_2_400_s_0_360 = 1.08e-04  mcm5m4p1_cc_w_2_400_s_0_360 = 1.00e-10  mcm5m4p1_cf_w_2_400_s_0_360 = 1.47e-11
+ mcm5m4p1_ca_w_2_400_s_0_450 = 1.08e-04  mcm5m4p1_cc_w_2_400_s_0_450 = 8.70e-11  mcm5m4p1_cf_w_2_400_s_0_450 = 1.82e-11
+ mcm5m4p1_ca_w_2_400_s_0_600 = 1.08e-04  mcm5m4p1_cc_w_2_400_s_0_600 = 7.03e-11  mcm5m4p1_cf_w_2_400_s_0_600 = 2.33e-11
+ mcm5m4p1_ca_w_2_400_s_0_800 = 1.08e-04  mcm5m4p1_cc_w_2_400_s_0_800 = 5.38e-11  mcm5m4p1_cf_w_2_400_s_0_800 = 2.94e-11
+ mcm5m4p1_ca_w_2_400_s_1_000 = 1.08e-04  mcm5m4p1_cc_w_2_400_s_1_000 = 4.21e-11  mcm5m4p1_cf_w_2_400_s_1_000 = 3.46e-11
+ mcm5m4p1_ca_w_2_400_s_1_200 = 1.08e-04  mcm5m4p1_cc_w_2_400_s_1_200 = 3.35e-11  mcm5m4p1_cf_w_2_400_s_1_200 = 3.89e-11
+ mcm5m4p1_ca_w_2_400_s_2_100 = 1.08e-04  mcm5m4p1_cc_w_2_400_s_2_100 = 1.41e-11  mcm5m4p1_cf_w_2_400_s_2_100 = 5.17e-11
+ mcm5m4p1_ca_w_2_400_s_3_300 = 1.08e-04  mcm5m4p1_cc_w_2_400_s_3_300 = 5.27e-12  mcm5m4p1_cf_w_2_400_s_3_300 = 5.93e-11
+ mcm5m4p1_ca_w_2_400_s_9_000 = 1.08e-04  mcm5m4p1_cc_w_2_400_s_9_000 = 1.30e-13  mcm5m4p1_cf_w_2_400_s_9_000 = 6.43e-11
+ mcm5m4l1_ca_w_0_300_s_0_300 = 1.10e-04  mcm5m4l1_cc_w_0_300_s_0_300 = 1.02e-10  mcm5m4l1_cf_w_0_300_s_0_300 = 1.24e-11
+ mcm5m4l1_ca_w_0_300_s_0_360 = 1.10e-04  mcm5m4l1_cc_w_0_300_s_0_360 = 9.22e-11  mcm5m4l1_cf_w_0_300_s_0_360 = 1.49e-11
+ mcm5m4l1_ca_w_0_300_s_0_450 = 1.10e-04  mcm5m4l1_cc_w_0_300_s_0_450 = 8.00e-11  mcm5m4l1_cf_w_0_300_s_0_450 = 1.84e-11
+ mcm5m4l1_ca_w_0_300_s_0_600 = 1.10e-04  mcm5m4l1_cc_w_0_300_s_0_600 = 6.39e-11  mcm5m4l1_cf_w_0_300_s_0_600 = 2.38e-11
+ mcm5m4l1_ca_w_0_300_s_0_800 = 1.10e-04  mcm5m4l1_cc_w_0_300_s_0_800 = 4.85e-11  mcm5m4l1_cf_w_0_300_s_0_800 = 2.98e-11
+ mcm5m4l1_ca_w_0_300_s_1_000 = 1.10e-04  mcm5m4l1_cc_w_0_300_s_1_000 = 3.74e-11  mcm5m4l1_cf_w_0_300_s_1_000 = 3.51e-11
+ mcm5m4l1_ca_w_0_300_s_1_200 = 1.10e-04  mcm5m4l1_cc_w_0_300_s_1_200 = 2.93e-11  mcm5m4l1_cf_w_0_300_s_1_200 = 3.94e-11
+ mcm5m4l1_ca_w_0_300_s_2_100 = 1.10e-04  mcm5m4l1_cc_w_0_300_s_2_100 = 1.14e-11  mcm5m4l1_cf_w_0_300_s_2_100 = 5.19e-11
+ mcm5m4l1_ca_w_0_300_s_3_300 = 1.10e-04  mcm5m4l1_cc_w_0_300_s_3_300 = 3.85e-12  mcm5m4l1_cf_w_0_300_s_3_300 = 5.86e-11
+ mcm5m4l1_ca_w_0_300_s_9_000 = 1.10e-04  mcm5m4l1_cc_w_0_300_s_9_000 = 6.50e-14  mcm5m4l1_cf_w_0_300_s_9_000 = 6.24e-11
+ mcm5m4l1_ca_w_2_400_s_0_300 = 1.10e-04  mcm5m4l1_cc_w_2_400_s_0_300 = 1.09e-10  mcm5m4l1_cf_w_2_400_s_0_300 = 1.24e-11
+ mcm5m4l1_ca_w_2_400_s_0_360 = 1.10e-04  mcm5m4l1_cc_w_2_400_s_0_360 = 9.90e-11  mcm5m4l1_cf_w_2_400_s_0_360 = 1.49e-11
+ mcm5m4l1_ca_w_2_400_s_0_450 = 1.10e-04  mcm5m4l1_cc_w_2_400_s_0_450 = 8.57e-11  mcm5m4l1_cf_w_2_400_s_0_450 = 1.85e-11
+ mcm5m4l1_ca_w_2_400_s_0_600 = 1.10e-04  mcm5m4l1_cc_w_2_400_s_0_600 = 6.91e-11  mcm5m4l1_cf_w_2_400_s_0_600 = 2.37e-11
+ mcm5m4l1_ca_w_2_400_s_0_800 = 1.10e-04  mcm5m4l1_cc_w_2_400_s_0_800 = 5.27e-11  mcm5m4l1_cf_w_2_400_s_0_800 = 2.99e-11
+ mcm5m4l1_ca_w_2_400_s_1_000 = 1.10e-04  mcm5m4l1_cc_w_2_400_s_1_000 = 4.07e-11  mcm5m4l1_cf_w_2_400_s_1_000 = 3.51e-11
+ mcm5m4l1_ca_w_2_400_s_1_200 = 1.10e-04  mcm5m4l1_cc_w_2_400_s_1_200 = 3.23e-11  mcm5m4l1_cf_w_2_400_s_1_200 = 3.96e-11
+ mcm5m4l1_ca_w_2_400_s_2_100 = 1.10e-04  mcm5m4l1_cc_w_2_400_s_2_100 = 1.31e-11  mcm5m4l1_cf_w_2_400_s_2_100 = 5.25e-11
+ mcm5m4l1_ca_w_2_400_s_3_300 = 1.10e-04  mcm5m4l1_cc_w_2_400_s_3_300 = 4.57e-12  mcm5m4l1_cf_w_2_400_s_3_300 = 5.99e-11
+ mcm5m4l1_ca_w_2_400_s_9_000 = 1.10e-04  mcm5m4l1_cc_w_2_400_s_9_000 = 9.00e-14  mcm5m4l1_cf_w_2_400_s_9_000 = 6.43e-11
+ mcm5m4m1_ca_w_0_300_s_0_300 = 1.14e-04  mcm5m4m1_cc_w_0_300_s_0_300 = 1.01e-10  mcm5m4m1_cf_w_0_300_s_0_300 = 1.29e-11
+ mcm5m4m1_ca_w_0_300_s_0_360 = 1.14e-04  mcm5m4m1_cc_w_0_300_s_0_360 = 9.11e-11  mcm5m4m1_cf_w_0_300_s_0_360 = 1.55e-11
+ mcm5m4m1_ca_w_0_300_s_0_450 = 1.14e-04  mcm5m4m1_cc_w_0_300_s_0_450 = 7.86e-11  mcm5m4m1_cf_w_0_300_s_0_450 = 1.92e-11
+ mcm5m4m1_ca_w_0_300_s_0_600 = 1.14e-04  mcm5m4m1_cc_w_0_300_s_0_600 = 6.26e-11  mcm5m4m1_cf_w_0_300_s_0_600 = 2.48e-11
+ mcm5m4m1_ca_w_0_300_s_0_800 = 1.14e-04  mcm5m4m1_cc_w_0_300_s_0_800 = 4.70e-11  mcm5m4m1_cf_w_0_300_s_0_800 = 3.12e-11
+ mcm5m4m1_ca_w_0_300_s_1_000 = 1.14e-04  mcm5m4m1_cc_w_0_300_s_1_000 = 3.58e-11  mcm5m4m1_cf_w_0_300_s_1_000 = 3.67e-11
+ mcm5m4m1_ca_w_0_300_s_1_200 = 1.14e-04  mcm5m4m1_cc_w_0_300_s_1_200 = 2.77e-11  mcm5m4m1_cf_w_0_300_s_1_200 = 4.11e-11
+ mcm5m4m1_ca_w_0_300_s_2_100 = 1.14e-04  mcm5m4m1_cc_w_0_300_s_2_100 = 1.00e-11  mcm5m4m1_cf_w_0_300_s_2_100 = 5.38e-11
+ mcm5m4m1_ca_w_0_300_s_3_300 = 1.14e-04  mcm5m4m1_cc_w_0_300_s_3_300 = 2.93e-12  mcm5m4m1_cf_w_0_300_s_3_300 = 6.02e-11
+ mcm5m4m1_ca_w_0_300_s_9_000 = 1.14e-04  mcm5m4m1_cc_w_0_300_s_9_000 = 6.00e-14  mcm5m4m1_cf_w_0_300_s_9_000 = 6.32e-11
+ mcm5m4m1_ca_w_2_400_s_0_300 = 1.14e-04  mcm5m4m1_cc_w_2_400_s_0_300 = 1.07e-10  mcm5m4m1_cf_w_2_400_s_0_300 = 1.29e-11
+ mcm5m4m1_ca_w_2_400_s_0_360 = 1.14e-04  mcm5m4m1_cc_w_2_400_s_0_360 = 9.64e-11  mcm5m4m1_cf_w_2_400_s_0_360 = 1.55e-11
+ mcm5m4m1_ca_w_2_400_s_0_450 = 1.14e-04  mcm5m4m1_cc_w_2_400_s_0_450 = 8.30e-11  mcm5m4m1_cf_w_2_400_s_0_450 = 1.92e-11
+ mcm5m4m1_ca_w_2_400_s_0_600 = 1.14e-04  mcm5m4m1_cc_w_2_400_s_0_600 = 6.64e-11  mcm5m4m1_cf_w_2_400_s_0_600 = 2.48e-11
+ mcm5m4m1_ca_w_2_400_s_0_800 = 1.14e-04  mcm5m4m1_cc_w_2_400_s_0_800 = 5.00e-11  mcm5m4m1_cf_w_2_400_s_0_800 = 3.12e-11
+ mcm5m4m1_ca_w_2_400_s_1_000 = 1.14e-04  mcm5m4m1_cc_w_2_400_s_1_000 = 3.82e-11  mcm5m4m1_cf_w_2_400_s_1_000 = 3.68e-11
+ mcm5m4m1_ca_w_2_400_s_1_200 = 1.14e-04  mcm5m4m1_cc_w_2_400_s_1_200 = 2.96e-11  mcm5m4m1_cf_w_2_400_s_1_200 = 4.13e-11
+ mcm5m4m1_ca_w_2_400_s_2_100 = 1.14e-04  mcm5m4m1_cc_w_2_400_s_2_100 = 1.10e-11  mcm5m4m1_cf_w_2_400_s_2_100 = 5.45e-11
+ mcm5m4m1_ca_w_2_400_s_3_300 = 1.14e-04  mcm5m4m1_cc_w_2_400_s_3_300 = 3.31e-12  mcm5m4m1_cf_w_2_400_s_3_300 = 6.14e-11
+ mcm5m4m1_ca_w_2_400_s_9_000 = 1.14e-04  mcm5m4m1_cc_w_2_400_s_9_000 = 6.50e-14  mcm5m4m1_cf_w_2_400_s_9_000 = 6.46e-11
+ mcm5m4m2_ca_w_0_300_s_0_300 = 1.20e-04  mcm5m4m2_cc_w_0_300_s_0_300 = 9.95e-11  mcm5m4m2_cf_w_0_300_s_0_300 = 1.38e-11
+ mcm5m4m2_ca_w_0_300_s_0_360 = 1.20e-04  mcm5m4m2_cc_w_0_300_s_0_360 = 8.94e-11  mcm5m4m2_cf_w_0_300_s_0_360 = 1.65e-11
+ mcm5m4m2_ca_w_0_300_s_0_450 = 1.20e-04  mcm5m4m2_cc_w_0_300_s_0_450 = 7.69e-11  mcm5m4m2_cf_w_0_300_s_0_450 = 2.05e-11
+ mcm5m4m2_ca_w_0_300_s_0_600 = 1.20e-04  mcm5m4m2_cc_w_0_300_s_0_600 = 6.07e-11  mcm5m4m2_cf_w_0_300_s_0_600 = 2.64e-11
+ mcm5m4m2_ca_w_0_300_s_0_800 = 1.20e-04  mcm5m4m2_cc_w_0_300_s_0_800 = 4.49e-11  mcm5m4m2_cf_w_0_300_s_0_800 = 3.33e-11
+ mcm5m4m2_ca_w_0_300_s_1_000 = 1.20e-04  mcm5m4m2_cc_w_0_300_s_1_000 = 3.36e-11  mcm5m4m2_cf_w_0_300_s_1_000 = 3.92e-11
+ mcm5m4m2_ca_w_0_300_s_1_200 = 1.20e-04  mcm5m4m2_cc_w_0_300_s_1_200 = 2.54e-11  mcm5m4m2_cf_w_0_300_s_1_200 = 4.40e-11
+ mcm5m4m2_ca_w_0_300_s_2_100 = 1.20e-04  mcm5m4m2_cc_w_0_300_s_2_100 = 8.15e-12  mcm5m4m2_cf_w_0_300_s_2_100 = 5.68e-11
+ mcm5m4m2_ca_w_0_300_s_3_300 = 1.20e-04  mcm5m4m2_cc_w_0_300_s_3_300 = 1.97e-12  mcm5m4m2_cf_w_0_300_s_3_300 = 6.26e-11
+ mcm5m4m2_ca_w_0_300_s_9_000 = 1.20e-04  mcm5m4m2_cc_w_0_300_s_9_000 = 4.00e-14  mcm5m4m2_cf_w_0_300_s_9_000 = 6.46e-11
+ mcm5m4m2_ca_w_2_400_s_0_300 = 1.20e-04  mcm5m4m2_cc_w_2_400_s_0_300 = 1.03e-10  mcm5m4m2_cf_w_2_400_s_0_300 = 1.38e-11
+ mcm5m4m2_ca_w_2_400_s_0_360 = 1.20e-04  mcm5m4m2_cc_w_2_400_s_0_360 = 9.30e-11  mcm5m4m2_cf_w_2_400_s_0_360 = 1.65e-11
+ mcm5m4m2_ca_w_2_400_s_0_450 = 1.20e-04  mcm5m4m2_cc_w_2_400_s_0_450 = 7.98e-11  mcm5m4m2_cf_w_2_400_s_0_450 = 2.05e-11
+ mcm5m4m2_ca_w_2_400_s_0_600 = 1.20e-04  mcm5m4m2_cc_w_2_400_s_0_600 = 6.30e-11  mcm5m4m2_cf_w_2_400_s_0_600 = 2.64e-11
+ mcm5m4m2_ca_w_2_400_s_0_800 = 1.20e-04  mcm5m4m2_cc_w_2_400_s_0_800 = 4.66e-11  mcm5m4m2_cf_w_2_400_s_0_800 = 3.34e-11
+ mcm5m4m2_ca_w_2_400_s_1_000 = 1.20e-04  mcm5m4m2_cc_w_2_400_s_1_000 = 3.49e-11  mcm5m4m2_cf_w_2_400_s_1_000 = 3.93e-11
+ mcm5m4m2_ca_w_2_400_s_1_200 = 1.20e-04  mcm5m4m2_cc_w_2_400_s_1_200 = 2.65e-11  mcm5m4m2_cf_w_2_400_s_1_200 = 4.41e-11
+ mcm5m4m2_ca_w_2_400_s_2_100 = 1.20e-04  mcm5m4m2_cc_w_2_400_s_2_100 = 8.60e-12  mcm5m4m2_cf_w_2_400_s_2_100 = 5.74e-11
+ mcm5m4m2_ca_w_2_400_s_3_300 = 1.20e-04  mcm5m4m2_cc_w_2_400_s_3_300 = 2.17e-12  mcm5m4m2_cf_w_2_400_s_3_300 = 6.34e-11
+ mcm5m4m2_ca_w_2_400_s_9_000 = 1.20e-04  mcm5m4m2_cc_w_2_400_s_9_000 = 1.50e-14  mcm5m4m2_cf_w_2_400_s_9_000 = 6.56e-11
+ mcm5m4m3_ca_w_0_300_s_0_300 = 2.38e-04  mcm5m4m3_cc_w_0_300_s_0_300 = 8.39e-11  mcm5m4m3_cf_w_0_300_s_0_300 = 2.68e-11
+ mcm5m4m3_ca_w_0_300_s_0_360 = 2.38e-04  mcm5m4m3_cc_w_0_300_s_0_360 = 7.37e-11  mcm5m4m3_cf_w_0_300_s_0_360 = 3.18e-11
+ mcm5m4m3_ca_w_0_300_s_0_450 = 2.38e-04  mcm5m4m3_cc_w_0_300_s_0_450 = 6.13e-11  mcm5m4m3_cf_w_0_300_s_0_450 = 3.87e-11
+ mcm5m4m3_ca_w_0_300_s_0_600 = 2.38e-04  mcm5m4m3_cc_w_0_300_s_0_600 = 4.49e-11  mcm5m4m3_cf_w_0_300_s_0_600 = 4.86e-11
+ mcm5m4m3_ca_w_0_300_s_0_800 = 2.38e-04  mcm5m4m3_cc_w_0_300_s_0_800 = 2.98e-11  mcm5m4m3_cf_w_0_300_s_0_800 = 5.89e-11
+ mcm5m4m3_ca_w_0_300_s_1_000 = 2.38e-04  mcm5m4m3_cc_w_0_300_s_1_000 = 1.94e-11  mcm5m4m3_cf_w_0_300_s_1_000 = 6.68e-11
+ mcm5m4m3_ca_w_0_300_s_1_200 = 2.38e-04  mcm5m4m3_cc_w_0_300_s_1_200 = 1.26e-11  mcm5m4m3_cf_w_0_300_s_1_200 = 7.23e-11
+ mcm5m4m3_ca_w_0_300_s_2_100 = 2.38e-04  mcm5m4m3_cc_w_0_300_s_2_100 = 2.00e-12  mcm5m4m3_cf_w_0_300_s_2_100 = 8.23e-11
+ mcm5m4m3_ca_w_0_300_s_3_300 = 2.38e-04  mcm5m4m3_cc_w_0_300_s_3_300 = 2.50e-13  mcm5m4m3_cf_w_0_300_s_3_300 = 8.45e-11
+ mcm5m4m3_ca_w_0_300_s_9_000 = 2.38e-04  mcm5m4m3_cc_w_0_300_s_9_000 = 5.00e-14  mcm5m4m3_cf_w_0_300_s_9_000 = 8.48e-11
+ mcm5m4m3_ca_w_2_400_s_0_300 = 2.38e-04  mcm5m4m3_cc_w_2_400_s_0_300 = 8.42e-11  mcm5m4m3_cf_w_2_400_s_0_300 = 2.67e-11
+ mcm5m4m3_ca_w_2_400_s_0_360 = 2.38e-04  mcm5m4m3_cc_w_2_400_s_0_360 = 7.42e-11  mcm5m4m3_cf_w_2_400_s_0_360 = 3.18e-11
+ mcm5m4m3_ca_w_2_400_s_0_450 = 2.38e-04  mcm5m4m3_cc_w_2_400_s_0_450 = 6.13e-11  mcm5m4m3_cf_w_2_400_s_0_450 = 3.87e-11
+ mcm5m4m3_ca_w_2_400_s_0_600 = 2.38e-04  mcm5m4m3_cc_w_2_400_s_0_600 = 4.51e-11  mcm5m4m3_cf_w_2_400_s_0_600 = 4.85e-11
+ mcm5m4m3_ca_w_2_400_s_0_800 = 2.38e-04  mcm5m4m3_cc_w_2_400_s_0_800 = 2.98e-11  mcm5m4m3_cf_w_2_400_s_0_800 = 5.90e-11
+ mcm5m4m3_ca_w_2_400_s_1_000 = 2.38e-04  mcm5m4m3_cc_w_2_400_s_1_000 = 1.94e-11  mcm5m4m3_cf_w_2_400_s_1_000 = 6.71e-11
+ mcm5m4m3_ca_w_2_400_s_1_200 = 2.38e-04  mcm5m4m3_cc_w_2_400_s_1_200 = 1.27e-11  mcm5m4m3_cf_w_2_400_s_1_200 = 7.26e-11
+ mcm5m4m3_ca_w_2_400_s_2_100 = 2.38e-04  mcm5m4m3_cc_w_2_400_s_2_100 = 1.95e-12  mcm5m4m3_cf_w_2_400_s_2_100 = 8.29e-11
+ mcm5m4m3_ca_w_2_400_s_3_300 = 2.38e-04  mcm5m4m3_cc_w_2_400_s_3_300 = 2.00e-13  mcm5m4m3_cf_w_2_400_s_3_300 = 8.47e-11
+ mcm5m4m3_ca_w_2_400_s_9_000 = 2.38e-04  mcm5m4m3_cc_w_2_400_s_9_000 = 0.00e+00  mcm5m4m3_cf_w_2_400_s_9_000 = 8.51e-11
+ mcrdlm4f_ca_w_0_300_s_0_300 = 1.55e-05  mcrdlm4f_cc_w_0_300_s_0_300 = 1.20e-10  mcrdlm4f_cf_w_0_300_s_0_300 = 2.04e-12
+ mcrdlm4f_ca_w_0_300_s_0_360 = 1.55e-05  mcrdlm4f_cc_w_0_300_s_0_360 = 1.11e-10  mcrdlm4f_cf_w_0_300_s_0_360 = 2.50e-12
+ mcrdlm4f_ca_w_0_300_s_0_450 = 1.55e-05  mcrdlm4f_cc_w_0_300_s_0_450 = 9.92e-11  mcrdlm4f_cf_w_0_300_s_0_450 = 3.22e-12
+ mcrdlm4f_ca_w_0_300_s_0_600 = 1.55e-05  mcrdlm4f_cc_w_0_300_s_0_600 = 8.49e-11  mcrdlm4f_cf_w_0_300_s_0_600 = 4.39e-12
+ mcrdlm4f_ca_w_0_300_s_0_800 = 1.55e-05  mcrdlm4f_cc_w_0_300_s_0_800 = 7.09e-11  mcrdlm4f_cf_w_0_300_s_0_800 = 5.75e-12
+ mcrdlm4f_ca_w_0_300_s_1_000 = 1.55e-05  mcrdlm4f_cc_w_0_300_s_1_000 = 6.07e-11  mcrdlm4f_cf_w_0_300_s_1_000 = 7.19e-12
+ mcrdlm4f_ca_w_0_300_s_1_200 = 1.55e-05  mcrdlm4f_cc_w_0_300_s_1_200 = 5.29e-11  mcrdlm4f_cf_w_0_300_s_1_200 = 8.58e-12
+ mcrdlm4f_ca_w_0_300_s_2_100 = 1.55e-05  mcrdlm4f_cc_w_0_300_s_2_100 = 3.31e-11  mcrdlm4f_cf_w_0_300_s_2_100 = 1.45e-11
+ mcrdlm4f_ca_w_0_300_s_3_300 = 1.55e-05  mcrdlm4f_cc_w_0_300_s_3_300 = 2.09e-11  mcrdlm4f_cf_w_0_300_s_3_300 = 2.04e-11
+ mcrdlm4f_ca_w_0_300_s_9_000 = 1.55e-05  mcrdlm4f_cc_w_0_300_s_9_000 = 3.40e-12  mcrdlm4f_cf_w_0_300_s_9_000 = 3.34e-11
+ mcrdlm4f_ca_w_2_400_s_0_300 = 1.55e-05  mcrdlm4f_cc_w_2_400_s_0_300 = 1.44e-10  mcrdlm4f_cf_w_2_400_s_0_300 = 2.08e-12
+ mcrdlm4f_ca_w_2_400_s_0_360 = 1.55e-05  mcrdlm4f_cc_w_2_400_s_0_360 = 1.34e-10  mcrdlm4f_cf_w_2_400_s_0_360 = 2.53e-12
+ mcrdlm4f_ca_w_2_400_s_0_450 = 1.55e-05  mcrdlm4f_cc_w_2_400_s_0_450 = 1.21e-10  mcrdlm4f_cf_w_2_400_s_0_450 = 3.21e-12
+ mcrdlm4f_ca_w_2_400_s_0_600 = 1.55e-05  mcrdlm4f_cc_w_2_400_s_0_600 = 1.04e-10  mcrdlm4f_cf_w_2_400_s_0_600 = 4.34e-12
+ mcrdlm4f_ca_w_2_400_s_0_800 = 1.55e-05  mcrdlm4f_cc_w_2_400_s_0_800 = 8.67e-11  mcrdlm4f_cf_w_2_400_s_0_800 = 5.81e-12
+ mcrdlm4f_ca_w_2_400_s_1_000 = 1.55e-05  mcrdlm4f_cc_w_2_400_s_1_000 = 7.43e-11  mcrdlm4f_cf_w_2_400_s_1_000 = 7.26e-12
+ mcrdlm4f_ca_w_2_400_s_1_200 = 1.55e-05  mcrdlm4f_cc_w_2_400_s_1_200 = 6.49e-11  mcrdlm4f_cf_w_2_400_s_1_200 = 8.67e-12
+ mcrdlm4f_ca_w_2_400_s_2_100 = 1.55e-05  mcrdlm4f_cc_w_2_400_s_2_100 = 4.11e-11  mcrdlm4f_cf_w_2_400_s_2_100 = 1.45e-11
+ mcrdlm4f_ca_w_2_400_s_3_300 = 1.55e-05  mcrdlm4f_cc_w_2_400_s_3_300 = 2.59e-11  mcrdlm4f_cf_w_2_400_s_3_300 = 2.11e-11
+ mcrdlm4f_ca_w_2_400_s_9_000 = 1.55e-05  mcrdlm4f_cc_w_2_400_s_9_000 = 4.36e-12  mcrdlm4f_cf_w_2_400_s_9_000 = 3.64e-11
+ mcrdlm4d_ca_w_0_300_s_0_300 = 1.63e-05  mcrdlm4d_cc_w_0_300_s_0_300 = 1.19e-10  mcrdlm4d_cf_w_0_300_s_0_300 = 2.14e-12
+ mcrdlm4d_ca_w_0_300_s_0_360 = 1.63e-05  mcrdlm4d_cc_w_0_300_s_0_360 = 1.11e-10  mcrdlm4d_cf_w_0_300_s_0_360 = 2.62e-12
+ mcrdlm4d_ca_w_0_300_s_0_450 = 1.63e-05  mcrdlm4d_cc_w_0_300_s_0_450 = 9.90e-11  mcrdlm4d_cf_w_0_300_s_0_450 = 3.37e-12
+ mcrdlm4d_ca_w_0_300_s_0_600 = 1.63e-05  mcrdlm4d_cc_w_0_300_s_0_600 = 8.47e-11  mcrdlm4d_cf_w_0_300_s_0_600 = 4.59e-12
+ mcrdlm4d_ca_w_0_300_s_0_800 = 1.63e-05  mcrdlm4d_cc_w_0_300_s_0_800 = 7.06e-11  mcrdlm4d_cf_w_0_300_s_0_800 = 6.01e-12
+ mcrdlm4d_ca_w_0_300_s_1_000 = 1.63e-05  mcrdlm4d_cc_w_0_300_s_1_000 = 6.03e-11  mcrdlm4d_cf_w_0_300_s_1_000 = 7.51e-12
+ mcrdlm4d_ca_w_0_300_s_1_200 = 1.63e-05  mcrdlm4d_cc_w_0_300_s_1_200 = 5.25e-11  mcrdlm4d_cf_w_0_300_s_1_200 = 8.97e-12
+ mcrdlm4d_ca_w_0_300_s_2_100 = 1.63e-05  mcrdlm4d_cc_w_0_300_s_2_100 = 3.27e-11  mcrdlm4d_cf_w_0_300_s_2_100 = 1.51e-11
+ mcrdlm4d_ca_w_0_300_s_3_300 = 1.63e-05  mcrdlm4d_cc_w_0_300_s_3_300 = 2.04e-11  mcrdlm4d_cf_w_0_300_s_3_300 = 2.11e-11
+ mcrdlm4d_ca_w_0_300_s_9_000 = 1.63e-05  mcrdlm4d_cc_w_0_300_s_9_000 = 3.17e-12  mcrdlm4d_cf_w_0_300_s_9_000 = 3.41e-11
+ mcrdlm4d_ca_w_2_400_s_0_300 = 1.63e-05  mcrdlm4d_cc_w_2_400_s_0_300 = 1.44e-10  mcrdlm4d_cf_w_2_400_s_0_300 = 2.18e-12
+ mcrdlm4d_ca_w_2_400_s_0_360 = 1.63e-05  mcrdlm4d_cc_w_2_400_s_0_360 = 1.34e-10  mcrdlm4d_cf_w_2_400_s_0_360 = 2.65e-12
+ mcrdlm4d_ca_w_2_400_s_0_450 = 1.63e-05  mcrdlm4d_cc_w_2_400_s_0_450 = 1.20e-10  mcrdlm4d_cf_w_2_400_s_0_450 = 3.36e-12
+ mcrdlm4d_ca_w_2_400_s_0_600 = 1.63e-05  mcrdlm4d_cc_w_2_400_s_0_600 = 1.03e-10  mcrdlm4d_cf_w_2_400_s_0_600 = 4.54e-12
+ mcrdlm4d_ca_w_2_400_s_0_800 = 1.63e-05  mcrdlm4d_cc_w_2_400_s_0_800 = 8.60e-11  mcrdlm4d_cf_w_2_400_s_0_800 = 6.08e-12
+ mcrdlm4d_ca_w_2_400_s_1_000 = 1.63e-05  mcrdlm4d_cc_w_2_400_s_1_000 = 7.37e-11  mcrdlm4d_cf_w_2_400_s_1_000 = 7.59e-12
+ mcrdlm4d_ca_w_2_400_s_1_200 = 1.63e-05  mcrdlm4d_cc_w_2_400_s_1_200 = 6.42e-11  mcrdlm4d_cf_w_2_400_s_1_200 = 9.05e-12
+ mcrdlm4d_ca_w_2_400_s_2_100 = 1.63e-05  mcrdlm4d_cc_w_2_400_s_2_100 = 4.04e-11  mcrdlm4d_cf_w_2_400_s_2_100 = 1.52e-11
+ mcrdlm4d_ca_w_2_400_s_3_300 = 1.63e-05  mcrdlm4d_cc_w_2_400_s_3_300 = 2.52e-11  mcrdlm4d_cf_w_2_400_s_3_300 = 2.19e-11
+ mcrdlm4d_ca_w_2_400_s_9_000 = 1.63e-05  mcrdlm4d_cc_w_2_400_s_9_000 = 4.11e-12  mcrdlm4d_cf_w_2_400_s_9_000 = 3.72e-11
+ mcrdlm4p1_ca_w_0_300_s_0_300 = 1.73e-05  mcrdlm4p1_cc_w_0_300_s_0_300 = 1.19e-10  mcrdlm4p1_cf_w_0_300_s_0_300 = 2.28e-12
+ mcrdlm4p1_ca_w_0_300_s_0_360 = 1.73e-05  mcrdlm4p1_cc_w_0_300_s_0_360 = 1.10e-10  mcrdlm4p1_cf_w_0_300_s_0_360 = 2.79e-12
+ mcrdlm4p1_ca_w_0_300_s_0_450 = 1.73e-05  mcrdlm4p1_cc_w_0_300_s_0_450 = 9.87e-11  mcrdlm4p1_cf_w_0_300_s_0_450 = 3.58e-12
+ mcrdlm4p1_ca_w_0_300_s_0_600 = 1.73e-05  mcrdlm4p1_cc_w_0_300_s_0_600 = 8.43e-11  mcrdlm4p1_cf_w_0_300_s_0_600 = 4.87e-12
+ mcrdlm4p1_ca_w_0_300_s_0_800 = 1.73e-05  mcrdlm4p1_cc_w_0_300_s_0_800 = 7.01e-11  mcrdlm4p1_cf_w_0_300_s_0_800 = 6.38e-12
+ mcrdlm4p1_ca_w_0_300_s_1_000 = 1.73e-05  mcrdlm4p1_cc_w_0_300_s_1_000 = 5.99e-11  mcrdlm4p1_cf_w_0_300_s_1_000 = 7.97e-12
+ mcrdlm4p1_ca_w_0_300_s_1_200 = 1.73e-05  mcrdlm4p1_cc_w_0_300_s_1_200 = 5.20e-11  mcrdlm4p1_cf_w_0_300_s_1_200 = 9.50e-12
+ mcrdlm4p1_ca_w_0_300_s_2_100 = 1.73e-05  mcrdlm4p1_cc_w_0_300_s_2_100 = 3.20e-11  mcrdlm4p1_cf_w_0_300_s_2_100 = 1.59e-11
+ mcrdlm4p1_ca_w_0_300_s_3_300 = 1.73e-05  mcrdlm4p1_cc_w_0_300_s_3_300 = 1.97e-11  mcrdlm4p1_cf_w_0_300_s_3_300 = 2.22e-11
+ mcrdlm4p1_ca_w_0_300_s_9_000 = 1.73e-05  mcrdlm4p1_cc_w_0_300_s_9_000 = 2.89e-12  mcrdlm4p1_cf_w_0_300_s_9_000 = 3.50e-11
+ mcrdlm4p1_ca_w_2_400_s_0_300 = 1.73e-05  mcrdlm4p1_cc_w_2_400_s_0_300 = 1.43e-10  mcrdlm4p1_cf_w_2_400_s_0_300 = 2.33e-12
+ mcrdlm4p1_ca_w_2_400_s_0_360 = 1.73e-05  mcrdlm4p1_cc_w_2_400_s_0_360 = 1.33e-10  mcrdlm4p1_cf_w_2_400_s_0_360 = 2.83e-12
+ mcrdlm4p1_ca_w_2_400_s_0_450 = 1.73e-05  mcrdlm4p1_cc_w_2_400_s_0_450 = 1.19e-10  mcrdlm4p1_cf_w_2_400_s_0_450 = 3.59e-12
+ mcrdlm4p1_ca_w_2_400_s_0_600 = 1.73e-05  mcrdlm4p1_cc_w_2_400_s_0_600 = 1.02e-10  mcrdlm4p1_cf_w_2_400_s_0_600 = 4.83e-12
+ mcrdlm4p1_ca_w_2_400_s_0_800 = 1.73e-05  mcrdlm4p1_cc_w_2_400_s_0_800 = 8.51e-11  mcrdlm4p1_cf_w_2_400_s_0_800 = 6.46e-12
+ mcrdlm4p1_ca_w_2_400_s_1_000 = 1.73e-05  mcrdlm4p1_cc_w_2_400_s_1_000 = 7.27e-11  mcrdlm4p1_cf_w_2_400_s_1_000 = 8.05e-12
+ mcrdlm4p1_ca_w_2_400_s_1_200 = 1.73e-05  mcrdlm4p1_cc_w_2_400_s_1_200 = 6.33e-11  mcrdlm4p1_cf_w_2_400_s_1_200 = 9.61e-12
+ mcrdlm4p1_ca_w_2_400_s_2_100 = 1.73e-05  mcrdlm4p1_cc_w_2_400_s_2_100 = 3.95e-11  mcrdlm4p1_cf_w_2_400_s_2_100 = 1.60e-11
+ mcrdlm4p1_ca_w_2_400_s_3_300 = 1.73e-05  mcrdlm4p1_cc_w_2_400_s_3_300 = 2.43e-11  mcrdlm4p1_cf_w_2_400_s_3_300 = 2.30e-11
+ mcrdlm4p1_ca_w_2_400_s_9_000 = 1.73e-05  mcrdlm4p1_cc_w_2_400_s_9_000 = 3.75e-12  mcrdlm4p1_cf_w_2_400_s_9_000 = 3.82e-11
+ mcrdlm4l1_ca_w_0_300_s_0_300 = 1.89e-05  mcrdlm4l1_cc_w_0_300_s_0_300 = 1.19e-10  mcrdlm4l1_cf_w_0_300_s_0_300 = 2.48e-12
+ mcrdlm4l1_ca_w_0_300_s_0_360 = 1.89e-05  mcrdlm4l1_cc_w_0_300_s_0_360 = 1.10e-10  mcrdlm4l1_cf_w_0_300_s_0_360 = 3.03e-12
+ mcrdlm4l1_ca_w_0_300_s_0_450 = 1.89e-05  mcrdlm4l1_cc_w_0_300_s_0_450 = 9.83e-11  mcrdlm4l1_cf_w_0_300_s_0_450 = 3.89e-12
+ mcrdlm4l1_ca_w_0_300_s_0_600 = 1.89e-05  mcrdlm4l1_cc_w_0_300_s_0_600 = 8.37e-11  mcrdlm4l1_cf_w_0_300_s_0_600 = 5.28e-12
+ mcrdlm4l1_ca_w_0_300_s_0_800 = 1.89e-05  mcrdlm4l1_cc_w_0_300_s_0_800 = 6.95e-11  mcrdlm4l1_cf_w_0_300_s_0_800 = 6.93e-12
+ mcrdlm4l1_ca_w_0_300_s_1_000 = 1.89e-05  mcrdlm4l1_cc_w_0_300_s_1_000 = 5.92e-11  mcrdlm4l1_cf_w_0_300_s_1_000 = 8.65e-12
+ mcrdlm4l1_ca_w_0_300_s_1_200 = 1.89e-05  mcrdlm4l1_cc_w_0_300_s_1_200 = 5.12e-11  mcrdlm4l1_cf_w_0_300_s_1_200 = 1.03e-11
+ mcrdlm4l1_ca_w_0_300_s_2_100 = 1.89e-05  mcrdlm4l1_cc_w_0_300_s_2_100 = 3.11e-11  mcrdlm4l1_cf_w_0_300_s_2_100 = 1.71e-11
+ mcrdlm4l1_ca_w_0_300_s_3_300 = 1.89e-05  mcrdlm4l1_cc_w_0_300_s_3_300 = 1.88e-11  mcrdlm4l1_cf_w_0_300_s_3_300 = 2.36e-11
+ mcrdlm4l1_ca_w_0_300_s_9_000 = 1.89e-05  mcrdlm4l1_cc_w_0_300_s_9_000 = 2.57e-12  mcrdlm4l1_cf_w_0_300_s_9_000 = 3.64e-11
+ mcrdlm4l1_ca_w_2_400_s_0_300 = 1.89e-05  mcrdlm4l1_cc_w_2_400_s_0_300 = 1.42e-10  mcrdlm4l1_cf_w_2_400_s_0_300 = 2.51e-12
+ mcrdlm4l1_ca_w_2_400_s_0_360 = 1.89e-05  mcrdlm4l1_cc_w_2_400_s_0_360 = 1.32e-10  mcrdlm4l1_cf_w_2_400_s_0_360 = 3.06e-12
+ mcrdlm4l1_ca_w_2_400_s_0_450 = 1.89e-05  mcrdlm4l1_cc_w_2_400_s_0_450 = 1.18e-10  mcrdlm4l1_cf_w_2_400_s_0_450 = 3.88e-12
+ mcrdlm4l1_ca_w_2_400_s_0_600 = 1.89e-05  mcrdlm4l1_cc_w_2_400_s_0_600 = 1.01e-10  mcrdlm4l1_cf_w_2_400_s_0_600 = 5.23e-12
+ mcrdlm4l1_ca_w_2_400_s_0_800 = 1.89e-05  mcrdlm4l1_cc_w_2_400_s_0_800 = 8.39e-11  mcrdlm4l1_cf_w_2_400_s_0_800 = 6.99e-12
+ mcrdlm4l1_ca_w_2_400_s_1_000 = 1.89e-05  mcrdlm4l1_cc_w_2_400_s_1_000 = 7.15e-11  mcrdlm4l1_cf_w_2_400_s_1_000 = 8.72e-12
+ mcrdlm4l1_ca_w_2_400_s_1_200 = 1.89e-05  mcrdlm4l1_cc_w_2_400_s_1_200 = 6.20e-11  mcrdlm4l1_cf_w_2_400_s_1_200 = 1.04e-11
+ mcrdlm4l1_ca_w_2_400_s_2_100 = 1.89e-05  mcrdlm4l1_cc_w_2_400_s_2_100 = 3.82e-11  mcrdlm4l1_cf_w_2_400_s_2_100 = 1.72e-11
+ mcrdlm4l1_ca_w_2_400_s_3_300 = 1.89e-05  mcrdlm4l1_cc_w_2_400_s_3_300 = 2.32e-11  mcrdlm4l1_cf_w_2_400_s_3_300 = 2.45e-11
+ mcrdlm4l1_ca_w_2_400_s_9_000 = 1.89e-05  mcrdlm4l1_cc_w_2_400_s_9_000 = 3.34e-12  mcrdlm4l1_cf_w_2_400_s_9_000 = 3.96e-11
+ mcrdlm4m1_ca_w_0_300_s_0_300 = 2.29e-05  mcrdlm4m1_cc_w_0_300_s_0_300 = 1.18e-10  mcrdlm4m1_cf_w_0_300_s_0_300 = 2.99e-12
+ mcrdlm4m1_ca_w_0_300_s_0_360 = 2.29e-05  mcrdlm4m1_cc_w_0_300_s_0_360 = 1.09e-10  mcrdlm4m1_cf_w_0_300_s_0_360 = 3.65e-12
+ mcrdlm4m1_ca_w_0_300_s_0_450 = 2.29e-05  mcrdlm4m1_cc_w_0_300_s_0_450 = 9.71e-11  mcrdlm4m1_cf_w_0_300_s_0_450 = 4.67e-12
+ mcrdlm4m1_ca_w_0_300_s_0_600 = 2.29e-05  mcrdlm4m1_cc_w_0_300_s_0_600 = 8.23e-11  mcrdlm4m1_cf_w_0_300_s_0_600 = 6.32e-12
+ mcrdlm4m1_ca_w_0_300_s_0_800 = 2.29e-05  mcrdlm4m1_cc_w_0_300_s_0_800 = 6.79e-11  mcrdlm4m1_cf_w_0_300_s_0_800 = 8.30e-12
+ mcrdlm4m1_ca_w_0_300_s_1_000 = 2.29e-05  mcrdlm4m1_cc_w_0_300_s_1_000 = 5.73e-11  mcrdlm4m1_cf_w_0_300_s_1_000 = 1.03e-11
+ mcrdlm4m1_ca_w_0_300_s_1_200 = 2.29e-05  mcrdlm4m1_cc_w_0_300_s_1_200 = 4.94e-11  mcrdlm4m1_cf_w_0_300_s_1_200 = 1.22e-11
+ mcrdlm4m1_ca_w_0_300_s_2_100 = 2.29e-05  mcrdlm4m1_cc_w_0_300_s_2_100 = 2.91e-11  mcrdlm4m1_cf_w_0_300_s_2_100 = 1.99e-11
+ mcrdlm4m1_ca_w_0_300_s_3_300 = 2.29e-05  mcrdlm4m1_cc_w_0_300_s_3_300 = 1.69e-11  mcrdlm4m1_cf_w_0_300_s_3_300 = 2.70e-11
+ mcrdlm4m1_ca_w_0_300_s_9_000 = 2.29e-05  mcrdlm4m1_cc_w_0_300_s_9_000 = 1.97e-12  mcrdlm4m1_cf_w_0_300_s_9_000 = 3.92e-11
+ mcrdlm4m1_ca_w_2_400_s_0_300 = 2.29e-05  mcrdlm4m1_cc_w_2_400_s_0_300 = 1.39e-10  mcrdlm4m1_cf_w_2_400_s_0_300 = 3.00e-12
+ mcrdlm4m1_ca_w_2_400_s_0_360 = 2.29e-05  mcrdlm4m1_cc_w_2_400_s_0_360 = 1.29e-10  mcrdlm4m1_cf_w_2_400_s_0_360 = 3.66e-12
+ mcrdlm4m1_ca_w_2_400_s_0_450 = 2.29e-05  mcrdlm4m1_cc_w_2_400_s_0_450 = 1.16e-10  mcrdlm4m1_cf_w_2_400_s_0_450 = 4.65e-12
+ mcrdlm4m1_ca_w_2_400_s_0_600 = 2.29e-05  mcrdlm4m1_cc_w_2_400_s_0_600 = 9.81e-11  mcrdlm4m1_cf_w_2_400_s_0_600 = 6.27e-12
+ mcrdlm4m1_ca_w_2_400_s_0_800 = 2.29e-05  mcrdlm4m1_cc_w_2_400_s_0_800 = 8.13e-11  mcrdlm4m1_cf_w_2_400_s_0_800 = 8.35e-12
+ mcrdlm4m1_ca_w_2_400_s_1_000 = 2.29e-05  mcrdlm4m1_cc_w_2_400_s_1_000 = 6.87e-11  mcrdlm4m1_cf_w_2_400_s_1_000 = 1.04e-11
+ mcrdlm4m1_ca_w_2_400_s_1_200 = 2.29e-05  mcrdlm4m1_cc_w_2_400_s_1_200 = 5.93e-11  mcrdlm4m1_cf_w_2_400_s_1_200 = 1.23e-11
+ mcrdlm4m1_ca_w_2_400_s_2_100 = 2.29e-05  mcrdlm4m1_cc_w_2_400_s_2_100 = 3.56e-11  mcrdlm4m1_cf_w_2_400_s_2_100 = 2.01e-11
+ mcrdlm4m1_ca_w_2_400_s_3_300 = 2.29e-05  mcrdlm4m1_cc_w_2_400_s_3_300 = 2.10e-11  mcrdlm4m1_cf_w_2_400_s_3_300 = 2.80e-11
+ mcrdlm4m1_ca_w_2_400_s_9_000 = 2.29e-05  mcrdlm4m1_cc_w_2_400_s_9_000 = 2.58e-12  mcrdlm4m1_cf_w_2_400_s_9_000 = 4.26e-11
+ mcrdlm4m2_ca_w_0_300_s_0_300 = 2.93e-05  mcrdlm4m2_cc_w_0_300_s_0_300 = 1.16e-10  mcrdlm4m2_cf_w_0_300_s_0_300 = 3.81e-12
+ mcrdlm4m2_ca_w_0_300_s_0_360 = 2.93e-05  mcrdlm4m2_cc_w_0_300_s_0_360 = 1.08e-10  mcrdlm4m2_cf_w_0_300_s_0_360 = 4.65e-12
+ mcrdlm4m2_ca_w_0_300_s_0_450 = 2.93e-05  mcrdlm4m2_cc_w_0_300_s_0_450 = 9.53e-11  mcrdlm4m2_cf_w_0_300_s_0_450 = 5.91e-12
+ mcrdlm4m2_ca_w_0_300_s_0_600 = 2.93e-05  mcrdlm4m2_cc_w_0_300_s_0_600 = 8.03e-11  mcrdlm4m2_cf_w_0_300_s_0_600 = 7.96e-12
+ mcrdlm4m2_ca_w_0_300_s_0_800 = 2.93e-05  mcrdlm4m2_cc_w_0_300_s_0_800 = 6.58e-11  mcrdlm4m2_cf_w_0_300_s_0_800 = 1.04e-11
+ mcrdlm4m2_ca_w_0_300_s_1_000 = 2.93e-05  mcrdlm4m2_cc_w_0_300_s_1_000 = 5.50e-11  mcrdlm4m2_cf_w_0_300_s_1_000 = 1.29e-11
+ mcrdlm4m2_ca_w_0_300_s_1_200 = 2.93e-05  mcrdlm4m2_cc_w_0_300_s_1_200 = 4.69e-11  mcrdlm4m2_cf_w_0_300_s_1_200 = 1.52e-11
+ mcrdlm4m2_ca_w_0_300_s_2_100 = 2.93e-05  mcrdlm4m2_cc_w_0_300_s_2_100 = 2.65e-11  mcrdlm4m2_cf_w_0_300_s_2_100 = 2.41e-11
+ mcrdlm4m2_ca_w_0_300_s_3_300 = 2.93e-05  mcrdlm4m2_cc_w_0_300_s_3_300 = 1.46e-11  mcrdlm4m2_cf_w_0_300_s_3_300 = 3.17e-11
+ mcrdlm4m2_ca_w_0_300_s_9_000 = 2.93e-05  mcrdlm4m2_cc_w_0_300_s_9_000 = 1.43e-12  mcrdlm4m2_cf_w_0_300_s_9_000 = 4.30e-11
+ mcrdlm4m2_ca_w_2_400_s_0_300 = 2.93e-05  mcrdlm4m2_cc_w_2_400_s_0_300 = 1.36e-10  mcrdlm4m2_cf_w_2_400_s_0_300 = 3.82e-12
+ mcrdlm4m2_ca_w_2_400_s_0_360 = 2.93e-05  mcrdlm4m2_cc_w_2_400_s_0_360 = 1.26e-10  mcrdlm4m2_cf_w_2_400_s_0_360 = 4.66e-12
+ mcrdlm4m2_ca_w_2_400_s_0_450 = 2.93e-05  mcrdlm4m2_cc_w_2_400_s_0_450 = 1.12e-10  mcrdlm4m2_cf_w_2_400_s_0_450 = 5.90e-12
+ mcrdlm4m2_ca_w_2_400_s_0_600 = 2.93e-05  mcrdlm4m2_cc_w_2_400_s_0_600 = 9.50e-11  mcrdlm4m2_cf_w_2_400_s_0_600 = 7.92e-12
+ mcrdlm4m2_ca_w_2_400_s_0_800 = 2.93e-05  mcrdlm4m2_cc_w_2_400_s_0_800 = 7.79e-11  mcrdlm4m2_cf_w_2_400_s_0_800 = 1.05e-11
+ mcrdlm4m2_ca_w_2_400_s_1_000 = 2.93e-05  mcrdlm4m2_cc_w_2_400_s_1_000 = 6.54e-11  mcrdlm4m2_cf_w_2_400_s_1_000 = 1.30e-11
+ mcrdlm4m2_ca_w_2_400_s_1_200 = 2.93e-05  mcrdlm4m2_cc_w_2_400_s_1_200 = 5.60e-11  mcrdlm4m2_cf_w_2_400_s_1_200 = 1.53e-11
+ mcrdlm4m2_ca_w_2_400_s_2_100 = 2.93e-05  mcrdlm4m2_cc_w_2_400_s_2_100 = 3.26e-11  mcrdlm4m2_cf_w_2_400_s_2_100 = 2.43e-11
+ mcrdlm4m2_ca_w_2_400_s_3_300 = 2.93e-05  mcrdlm4m2_cc_w_2_400_s_3_300 = 1.84e-11  mcrdlm4m2_cf_w_2_400_s_3_300 = 3.28e-11
+ mcrdlm4m2_ca_w_2_400_s_9_000 = 2.93e-05  mcrdlm4m2_cc_w_2_400_s_9_000 = 1.97e-12  mcrdlm4m2_cf_w_2_400_s_9_000 = 4.66e-11
+ mcrdlm4m3_ca_w_0_300_s_0_300 = 1.47e-04  mcrdlm4m3_cc_w_0_300_s_0_300 = 1.01e-10  mcrdlm4m3_cf_w_0_300_s_0_300 = 1.68e-11
+ mcrdlm4m3_ca_w_0_300_s_0_360 = 1.47e-04  mcrdlm4m3_cc_w_0_300_s_0_360 = 9.17e-11  mcrdlm4m3_cf_w_0_300_s_0_360 = 1.99e-11
+ mcrdlm4m3_ca_w_0_300_s_0_450 = 1.47e-04  mcrdlm4m3_cc_w_0_300_s_0_450 = 7.94e-11  mcrdlm4m3_cf_w_0_300_s_0_450 = 2.41e-11
+ mcrdlm4m3_ca_w_0_300_s_0_600 = 1.47e-04  mcrdlm4m3_cc_w_0_300_s_0_600 = 6.44e-11  mcrdlm4m3_cf_w_0_300_s_0_600 = 3.02e-11
+ mcrdlm4m3_ca_w_0_300_s_0_800 = 1.47e-04  mcrdlm4m3_cc_w_0_300_s_0_800 = 5.03e-11  mcrdlm4m3_cf_w_0_300_s_0_800 = 3.65e-11
+ mcrdlm4m3_ca_w_0_300_s_1_000 = 1.47e-04  mcrdlm4m3_cc_w_0_300_s_1_000 = 3.99e-11  mcrdlm4m3_cf_w_0_300_s_1_000 = 4.18e-11
+ mcrdlm4m3_ca_w_0_300_s_1_200 = 1.47e-04  mcrdlm4m3_cc_w_0_300_s_1_200 = 3.25e-11  mcrdlm4m3_cf_w_0_300_s_1_200 = 4.60e-11
+ mcrdlm4m3_ca_w_0_300_s_2_100 = 1.47e-04  mcrdlm4m3_cc_w_0_300_s_2_100 = 1.52e-11  mcrdlm4m3_cf_w_0_300_s_2_100 = 5.83e-11
+ mcrdlm4m3_ca_w_0_300_s_3_300 = 1.47e-04  mcrdlm4m3_cc_w_0_300_s_3_300 = 7.10e-12  mcrdlm4m3_cf_w_0_300_s_3_300 = 6.54e-11
+ mcrdlm4m3_ca_w_0_300_s_9_000 = 1.47e-04  mcrdlm4m3_cc_w_0_300_s_9_000 = 4.85e-13  mcrdlm4m3_cf_w_0_300_s_9_000 = 7.17e-11
+ mcrdlm4m3_ca_w_2_400_s_0_300 = 1.47e-04  mcrdlm4m3_cc_w_2_400_s_0_300 = 1.16e-10  mcrdlm4m3_cf_w_2_400_s_0_300 = 1.68e-11
+ mcrdlm4m3_ca_w_2_400_s_0_360 = 1.47e-04  mcrdlm4m3_cc_w_2_400_s_0_360 = 1.06e-10  mcrdlm4m3_cf_w_2_400_s_0_360 = 1.99e-11
+ mcrdlm4m3_ca_w_2_400_s_0_450 = 1.47e-04  mcrdlm4m3_cc_w_2_400_s_0_450 = 9.35e-11  mcrdlm4m3_cf_w_2_400_s_0_450 = 2.41e-11
+ mcrdlm4m3_ca_w_2_400_s_0_600 = 1.47e-04  mcrdlm4m3_cc_w_2_400_s_0_600 = 7.67e-11  mcrdlm4m3_cf_w_2_400_s_0_600 = 3.01e-11
+ mcrdlm4m3_ca_w_2_400_s_0_800 = 1.47e-04  mcrdlm4m3_cc_w_2_400_s_0_800 = 6.09e-11  mcrdlm4m3_cf_w_2_400_s_0_800 = 3.66e-11
+ mcrdlm4m3_ca_w_2_400_s_1_000 = 1.47e-04  mcrdlm4m3_cc_w_2_400_s_1_000 = 4.94e-11  mcrdlm4m3_cf_w_2_400_s_1_000 = 4.19e-11
+ mcrdlm4m3_ca_w_2_400_s_1_200 = 1.47e-04  mcrdlm4m3_cc_w_2_400_s_1_200 = 4.09e-11  mcrdlm4m3_cf_w_2_400_s_1_200 = 4.62e-11
+ mcrdlm4m3_ca_w_2_400_s_2_100 = 1.47e-04  mcrdlm4m3_cc_w_2_400_s_2_100 = 2.11e-11  mcrdlm4m3_cf_w_2_400_s_2_100 = 5.89e-11
+ mcrdlm4m3_ca_w_2_400_s_3_300 = 1.47e-04  mcrdlm4m3_cc_w_2_400_s_3_300 = 1.05e-11  mcrdlm4m3_cf_w_2_400_s_3_300 = 6.76e-11
+ mcrdlm4m3_ca_w_2_400_s_9_000 = 1.47e-04  mcrdlm4m3_cc_w_2_400_s_9_000 = 7.15e-13  mcrdlm4m3_cf_w_2_400_s_9_000 = 7.68e-11
+ mcrdlm5f_ca_w_1_600_s_1_600 = 1.53e-05  mcrdlm5f_cc_w_1_600_s_1_600 = 7.56e-11  mcrdlm5f_cf_w_1_600_s_1_600 = 1.11e-11
+ mcrdlm5f_ca_w_1_600_s_1_700 = 1.53e-05  mcrdlm5f_cc_w_1_600_s_1_700 = 7.09e-11  mcrdlm5f_cf_w_1_600_s_1_700 = 1.17e-11
+ mcrdlm5f_ca_w_1_600_s_1_900 = 1.53e-05  mcrdlm5f_cc_w_1_600_s_1_900 = 6.31e-11  mcrdlm5f_cf_w_1_600_s_1_900 = 1.31e-11
+ mcrdlm5f_ca_w_1_600_s_2_000 = 1.53e-05  mcrdlm5f_cc_w_1_600_s_2_000 = 5.98e-11  mcrdlm5f_cf_w_1_600_s_2_000 = 1.37e-11
+ mcrdlm5f_ca_w_1_600_s_2_400 = 1.53e-05  mcrdlm5f_cc_w_1_600_s_2_400 = 4.91e-11  mcrdlm5f_cf_w_1_600_s_2_400 = 1.63e-11
+ mcrdlm5f_ca_w_1_600_s_2_800 = 1.53e-05  mcrdlm5f_cc_w_1_600_s_2_800 = 4.12e-11  mcrdlm5f_cf_w_1_600_s_2_800 = 1.87e-11
+ mcrdlm5f_ca_w_1_600_s_3_200 = 1.53e-05  mcrdlm5f_cc_w_1_600_s_3_200 = 3.51e-11  mcrdlm5f_cf_w_1_600_s_3_200 = 2.10e-11
+ mcrdlm5f_ca_w_1_600_s_4_800 = 1.53e-05  mcrdlm5f_cc_w_1_600_s_4_800 = 2.01e-11  mcrdlm5f_cf_w_1_600_s_4_800 = 2.86e-11
+ mcrdlm5f_ca_w_1_600_s_10_000 = 1.53e-05  mcrdlm5f_cc_w_1_600_s_10_000 = 4.11e-12  mcrdlm5f_cf_w_1_600_s_10_000 = 4.07e-11
+ mcrdlm5f_ca_w_1_600_s_12_000 = 1.53e-05  mcrdlm5f_cc_w_1_600_s_12_000 = 2.29e-12  mcrdlm5f_cf_w_1_600_s_12_000 = 4.25e-11
+ mcrdlm5f_ca_w_4_000_s_1_600 = 1.53e-05  mcrdlm5f_cc_w_4_000_s_1_600 = 7.82e-11  mcrdlm5f_cf_w_4_000_s_1_600 = 1.11e-11
+ mcrdlm5f_ca_w_4_000_s_1_700 = 1.53e-05  mcrdlm5f_cc_w_4_000_s_1_700 = 7.33e-11  mcrdlm5f_cf_w_4_000_s_1_700 = 1.17e-11
+ mcrdlm5f_ca_w_4_000_s_1_900 = 1.53e-05  mcrdlm5f_cc_w_4_000_s_1_900 = 6.52e-11  mcrdlm5f_cf_w_4_000_s_1_900 = 1.31e-11
+ mcrdlm5f_ca_w_4_000_s_2_000 = 1.53e-05  mcrdlm5f_cc_w_4_000_s_2_000 = 6.18e-11  mcrdlm5f_cf_w_4_000_s_2_000 = 1.37e-11
+ mcrdlm5f_ca_w_4_000_s_2_400 = 1.53e-05  mcrdlm5f_cc_w_4_000_s_2_400 = 5.07e-11  mcrdlm5f_cf_w_4_000_s_2_400 = 1.63e-11
+ mcrdlm5f_ca_w_4_000_s_2_800 = 1.53e-05  mcrdlm5f_cc_w_4_000_s_2_800 = 4.26e-11  mcrdlm5f_cf_w_4_000_s_2_800 = 1.87e-11
+ mcrdlm5f_ca_w_4_000_s_3_200 = 1.53e-05  mcrdlm5f_cc_w_4_000_s_3_200 = 3.63e-11  mcrdlm5f_cf_w_4_000_s_3_200 = 2.10e-11
+ mcrdlm5f_ca_w_4_000_s_4_800 = 1.53e-05  mcrdlm5f_cc_w_4_000_s_4_800 = 2.08e-11  mcrdlm5f_cf_w_4_000_s_4_800 = 2.87e-11
+ mcrdlm5f_ca_w_4_000_s_10_000 = 1.53e-05  mcrdlm5f_cc_w_4_000_s_10_000 = 4.30e-12  mcrdlm5f_cf_w_4_000_s_10_000 = 4.13e-11
+ mcrdlm5f_ca_w_4_000_s_12_000 = 1.53e-05  mcrdlm5f_cc_w_4_000_s_12_000 = 2.40e-12  mcrdlm5f_cf_w_4_000_s_12_000 = 4.31e-11
+ mcrdlm5d_ca_w_1_600_s_1_600 = 1.57e-05  mcrdlm5d_cc_w_1_600_s_1_600 = 7.51e-11  mcrdlm5d_cf_w_1_600_s_1_600 = 1.13e-11
+ mcrdlm5d_ca_w_1_600_s_1_700 = 1.57e-05  mcrdlm5d_cc_w_1_600_s_1_700 = 7.05e-11  mcrdlm5d_cf_w_1_600_s_1_700 = 1.20e-11
+ mcrdlm5d_ca_w_1_600_s_1_900 = 1.57e-05  mcrdlm5d_cc_w_1_600_s_1_900 = 6.26e-11  mcrdlm5d_cf_w_1_600_s_1_900 = 1.34e-11
+ mcrdlm5d_ca_w_1_600_s_2_000 = 1.57e-05  mcrdlm5d_cc_w_1_600_s_2_000 = 5.94e-11  mcrdlm5d_cf_w_1_600_s_2_000 = 1.41e-11
+ mcrdlm5d_ca_w_1_600_s_2_400 = 1.57e-05  mcrdlm5d_cc_w_1_600_s_2_400 = 4.85e-11  mcrdlm5d_cf_w_1_600_s_2_400 = 1.66e-11
+ mcrdlm5d_ca_w_1_600_s_2_800 = 1.57e-05  mcrdlm5d_cc_w_1_600_s_2_800 = 4.07e-11  mcrdlm5d_cf_w_1_600_s_2_800 = 1.91e-11
+ mcrdlm5d_ca_w_1_600_s_3_200 = 1.57e-05  mcrdlm5d_cc_w_1_600_s_3_200 = 3.47e-11  mcrdlm5d_cf_w_1_600_s_3_200 = 2.14e-11
+ mcrdlm5d_ca_w_1_600_s_4_800 = 1.57e-05  mcrdlm5d_cc_w_1_600_s_4_800 = 1.97e-11  mcrdlm5d_cf_w_1_600_s_4_800 = 2.91e-11
+ mcrdlm5d_ca_w_1_600_s_10_000 = 1.57e-05  mcrdlm5d_cc_w_1_600_s_10_000 = 3.88e-12  mcrdlm5d_cf_w_1_600_s_10_000 = 4.13e-11
+ mcrdlm5d_ca_w_1_600_s_12_000 = 1.57e-05  mcrdlm5d_cc_w_1_600_s_12_000 = 2.12e-12  mcrdlm5d_cf_w_1_600_s_12_000 = 4.29e-11
+ mcrdlm5d_ca_w_4_000_s_1_600 = 1.57e-05  mcrdlm5d_cc_w_4_000_s_1_600 = 7.77e-11  mcrdlm5d_cf_w_4_000_s_1_600 = 1.13e-11
+ mcrdlm5d_ca_w_4_000_s_1_700 = 1.57e-05  mcrdlm5d_cc_w_4_000_s_1_700 = 7.28e-11  mcrdlm5d_cf_w_4_000_s_1_700 = 1.20e-11
+ mcrdlm5d_ca_w_4_000_s_1_900 = 1.57e-05  mcrdlm5d_cc_w_4_000_s_1_900 = 6.47e-11  mcrdlm5d_cf_w_4_000_s_1_900 = 1.34e-11
+ mcrdlm5d_ca_w_4_000_s_2_000 = 1.57e-05  mcrdlm5d_cc_w_4_000_s_2_000 = 6.13e-11  mcrdlm5d_cf_w_4_000_s_2_000 = 1.41e-11
+ mcrdlm5d_ca_w_4_000_s_2_400 = 1.57e-05  mcrdlm5d_cc_w_4_000_s_2_400 = 5.01e-11  mcrdlm5d_cf_w_4_000_s_2_400 = 1.67e-11
+ mcrdlm5d_ca_w_4_000_s_2_800 = 1.57e-05  mcrdlm5d_cc_w_4_000_s_2_800 = 4.20e-11  mcrdlm5d_cf_w_4_000_s_2_800 = 1.92e-11
+ mcrdlm5d_ca_w_4_000_s_3_200 = 1.57e-05  mcrdlm5d_cc_w_4_000_s_3_200 = 3.58e-11  mcrdlm5d_cf_w_4_000_s_3_200 = 2.15e-11
+ mcrdlm5d_ca_w_4_000_s_4_800 = 1.57e-05  mcrdlm5d_cc_w_4_000_s_4_800 = 2.04e-11  mcrdlm5d_cf_w_4_000_s_4_800 = 2.93e-11
+ mcrdlm5d_ca_w_4_000_s_10_000 = 1.57e-05  mcrdlm5d_cc_w_4_000_s_10_000 = 4.07e-12  mcrdlm5d_cf_w_4_000_s_10_000 = 4.18e-11
+ mcrdlm5d_ca_w_4_000_s_12_000 = 1.57e-05  mcrdlm5d_cc_w_4_000_s_12_000 = 2.24e-12  mcrdlm5d_cf_w_4_000_s_12_000 = 4.35e-11
+ mcrdlm5p1_ca_w_1_600_s_1_600 = 1.62e-05  mcrdlm5p1_cc_w_1_600_s_1_600 = 7.46e-11  mcrdlm5p1_cf_w_1_600_s_1_600 = 1.17e-11
+ mcrdlm5p1_ca_w_1_600_s_1_700 = 1.62e-05  mcrdlm5p1_cc_w_1_600_s_1_700 = 7.00e-11  mcrdlm5p1_cf_w_1_600_s_1_700 = 1.24e-11
+ mcrdlm5p1_ca_w_1_600_s_1_900 = 1.62e-05  mcrdlm5p1_cc_w_1_600_s_1_900 = 6.20e-11  mcrdlm5p1_cf_w_1_600_s_1_900 = 1.38e-11
+ mcrdlm5p1_ca_w_1_600_s_2_000 = 1.62e-05  mcrdlm5p1_cc_w_1_600_s_2_000 = 5.87e-11  mcrdlm5p1_cf_w_1_600_s_2_000 = 1.45e-11
+ mcrdlm5p1_ca_w_1_600_s_2_400 = 1.62e-05  mcrdlm5p1_cc_w_1_600_s_2_400 = 4.80e-11  mcrdlm5p1_cf_w_1_600_s_2_400 = 1.72e-11
+ mcrdlm5p1_ca_w_1_600_s_2_800 = 1.62e-05  mcrdlm5p1_cc_w_1_600_s_2_800 = 4.01e-11  mcrdlm5p1_cf_w_1_600_s_2_800 = 1.97e-11
+ mcrdlm5p1_ca_w_1_600_s_3_200 = 1.62e-05  mcrdlm5p1_cc_w_1_600_s_3_200 = 3.41e-11  mcrdlm5p1_cf_w_1_600_s_3_200 = 2.21e-11
+ mcrdlm5p1_ca_w_1_600_s_4_800 = 1.62e-05  mcrdlm5p1_cc_w_1_600_s_4_800 = 1.91e-11  mcrdlm5p1_cf_w_1_600_s_4_800 = 2.99e-11
+ mcrdlm5p1_ca_w_1_600_s_10_000 = 1.62e-05  mcrdlm5p1_cc_w_1_600_s_10_000 = 3.59e-12  mcrdlm5p1_cf_w_1_600_s_10_000 = 4.20e-11
+ mcrdlm5p1_ca_w_1_600_s_12_000 = 1.62e-05  mcrdlm5p1_cc_w_1_600_s_12_000 = 1.92e-12  mcrdlm5p1_cf_w_1_600_s_12_000 = 4.36e-11
+ mcrdlm5p1_ca_w_4_000_s_1_600 = 1.62e-05  mcrdlm5p1_cc_w_4_000_s_1_600 = 7.70e-11  mcrdlm5p1_cf_w_4_000_s_1_600 = 1.17e-11
+ mcrdlm5p1_ca_w_4_000_s_1_700 = 1.62e-05  mcrdlm5p1_cc_w_4_000_s_1_700 = 7.21e-11  mcrdlm5p1_cf_w_4_000_s_1_700 = 1.24e-11
+ mcrdlm5p1_ca_w_4_000_s_1_900 = 1.62e-05  mcrdlm5p1_cc_w_4_000_s_1_900 = 6.40e-11  mcrdlm5p1_cf_w_4_000_s_1_900 = 1.38e-11
+ mcrdlm5p1_ca_w_4_000_s_2_000 = 1.62e-05  mcrdlm5p1_cc_w_4_000_s_2_000 = 6.06e-11  mcrdlm5p1_cf_w_4_000_s_2_000 = 1.45e-11
+ mcrdlm5p1_ca_w_4_000_s_2_400 = 1.62e-05  mcrdlm5p1_cc_w_4_000_s_2_400 = 4.95e-11  mcrdlm5p1_cf_w_4_000_s_2_400 = 1.72e-11
+ mcrdlm5p1_ca_w_4_000_s_2_800 = 1.62e-05  mcrdlm5p1_cc_w_4_000_s_2_800 = 4.13e-11  mcrdlm5p1_cf_w_4_000_s_2_800 = 1.97e-11
+ mcrdlm5p1_ca_w_4_000_s_3_200 = 1.62e-05  mcrdlm5p1_cc_w_4_000_s_3_200 = 3.51e-11  mcrdlm5p1_cf_w_4_000_s_3_200 = 2.21e-11
+ mcrdlm5p1_ca_w_4_000_s_4_800 = 1.62e-05  mcrdlm5p1_cc_w_4_000_s_4_800 = 1.97e-11  mcrdlm5p1_cf_w_4_000_s_4_800 = 3.01e-11
+ mcrdlm5p1_ca_w_4_000_s_10_000 = 1.62e-05  mcrdlm5p1_cc_w_4_000_s_10_000 = 3.77e-12  mcrdlm5p1_cf_w_4_000_s_10_000 = 4.25e-11
+ mcrdlm5p1_ca_w_4_000_s_12_000 = 1.62e-05  mcrdlm5p1_cc_w_4_000_s_12_000 = 2.02e-12  mcrdlm5p1_cf_w_4_000_s_12_000 = 4.41e-11
+ mcrdlm5l1_ca_w_1_600_s_1_600 = 1.69e-05  mcrdlm5l1_cc_w_1_600_s_1_600 = 7.41e-11  mcrdlm5l1_cf_w_1_600_s_1_600 = 1.22e-11
+ mcrdlm5l1_ca_w_1_600_s_1_700 = 1.69e-05  mcrdlm5l1_cc_w_1_600_s_1_700 = 6.92e-11  mcrdlm5l1_cf_w_1_600_s_1_700 = 1.30e-11
+ mcrdlm5l1_ca_w_1_600_s_1_900 = 1.69e-05  mcrdlm5l1_cc_w_1_600_s_1_900 = 6.13e-11  mcrdlm5l1_cf_w_1_600_s_1_900 = 1.44e-11
+ mcrdlm5l1_ca_w_1_600_s_2_000 = 1.69e-05  mcrdlm5l1_cc_w_1_600_s_2_000 = 5.80e-11  mcrdlm5l1_cf_w_1_600_s_2_000 = 1.51e-11
+ mcrdlm5l1_ca_w_1_600_s_2_400 = 1.69e-05  mcrdlm5l1_cc_w_1_600_s_2_400 = 4.71e-11  mcrdlm5l1_cf_w_1_600_s_2_400 = 1.79e-11
+ mcrdlm5l1_ca_w_1_600_s_2_800 = 1.69e-05  mcrdlm5l1_cc_w_1_600_s_2_800 = 3.94e-11  mcrdlm5l1_cf_w_1_600_s_2_800 = 2.05e-11
+ mcrdlm5l1_ca_w_1_600_s_3_200 = 1.69e-05  mcrdlm5l1_cc_w_1_600_s_3_200 = 3.33e-11  mcrdlm5l1_cf_w_1_600_s_3_200 = 2.30e-11
+ mcrdlm5l1_ca_w_1_600_s_4_800 = 1.69e-05  mcrdlm5l1_cc_w_1_600_s_4_800 = 1.84e-11  mcrdlm5l1_cf_w_1_600_s_4_800 = 3.10e-11
+ mcrdlm5l1_ca_w_1_600_s_10_000 = 1.69e-05  mcrdlm5l1_cc_w_1_600_s_10_000 = 3.26e-12  mcrdlm5l1_cf_w_1_600_s_10_000 = 4.29e-11
+ mcrdlm5l1_ca_w_1_600_s_12_000 = 1.69e-05  mcrdlm5l1_cc_w_1_600_s_12_000 = 1.71e-12  mcrdlm5l1_cf_w_1_600_s_12_000 = 4.44e-11
+ mcrdlm5l1_ca_w_4_000_s_1_600 = 1.69e-05  mcrdlm5l1_cc_w_4_000_s_1_600 = 7.62e-11  mcrdlm5l1_cf_w_4_000_s_1_600 = 1.22e-11
+ mcrdlm5l1_ca_w_4_000_s_1_700 = 1.69e-05  mcrdlm5l1_cc_w_4_000_s_1_700 = 7.12e-11  mcrdlm5l1_cf_w_4_000_s_1_700 = 1.30e-11
+ mcrdlm5l1_ca_w_4_000_s_1_900 = 1.69e-05  mcrdlm5l1_cc_w_4_000_s_1_900 = 6.31e-11  mcrdlm5l1_cf_w_4_000_s_1_900 = 1.44e-11
+ mcrdlm5l1_ca_w_4_000_s_2_000 = 1.69e-05  mcrdlm5l1_cc_w_4_000_s_2_000 = 5.97e-11  mcrdlm5l1_cf_w_4_000_s_2_000 = 1.52e-11
+ mcrdlm5l1_ca_w_4_000_s_2_400 = 1.69e-05  mcrdlm5l1_cc_w_4_000_s_2_400 = 4.85e-11  mcrdlm5l1_cf_w_4_000_s_2_400 = 1.79e-11
+ mcrdlm5l1_ca_w_4_000_s_2_800 = 1.69e-05  mcrdlm5l1_cc_w_4_000_s_2_800 = 4.04e-11  mcrdlm5l1_cf_w_4_000_s_2_800 = 2.06e-11
+ mcrdlm5l1_ca_w_4_000_s_3_200 = 1.69e-05  mcrdlm5l1_cc_w_4_000_s_3_200 = 3.42e-11  mcrdlm5l1_cf_w_4_000_s_3_200 = 2.30e-11
+ mcrdlm5l1_ca_w_4_000_s_4_800 = 1.69e-05  mcrdlm5l1_cc_w_4_000_s_4_800 = 1.90e-11  mcrdlm5l1_cf_w_4_000_s_4_800 = 3.12e-11
+ mcrdlm5l1_ca_w_4_000_s_10_000 = 1.69e-05  mcrdlm5l1_cc_w_4_000_s_10_000 = 3.38e-12  mcrdlm5l1_cf_w_4_000_s_10_000 = 4.34e-11
+ mcrdlm5l1_ca_w_4_000_s_12_000 = 1.69e-05  mcrdlm5l1_cc_w_4_000_s_12_000 = 1.81e-12  mcrdlm5l1_cf_w_4_000_s_12_000 = 4.50e-11
+ mcrdlm5m1_ca_w_1_600_s_1_600 = 1.86e-05  mcrdlm5m1_cc_w_1_600_s_1_600 = 7.26e-11  mcrdlm5m1_cf_w_1_600_s_1_600 = 1.34e-11
+ mcrdlm5m1_ca_w_1_600_s_1_700 = 1.86e-05  mcrdlm5m1_cc_w_1_600_s_1_700 = 6.78e-11  mcrdlm5m1_cf_w_1_600_s_1_700 = 1.41e-11
+ mcrdlm5m1_ca_w_1_600_s_1_900 = 1.86e-05  mcrdlm5m1_cc_w_1_600_s_1_900 = 5.98e-11  mcrdlm5m1_cf_w_1_600_s_1_900 = 1.57e-11
+ mcrdlm5m1_ca_w_1_600_s_2_000 = 1.86e-05  mcrdlm5m1_cc_w_1_600_s_2_000 = 5.65e-11  mcrdlm5m1_cf_w_1_600_s_2_000 = 1.65e-11
+ mcrdlm5m1_ca_w_1_600_s_2_400 = 1.86e-05  mcrdlm5m1_cc_w_1_600_s_2_400 = 4.56e-11  mcrdlm5m1_cf_w_1_600_s_2_400 = 1.95e-11
+ mcrdlm5m1_ca_w_1_600_s_2_800 = 1.86e-05  mcrdlm5m1_cc_w_1_600_s_2_800 = 3.78e-11  mcrdlm5m1_cf_w_1_600_s_2_800 = 2.23e-11
+ mcrdlm5m1_ca_w_1_600_s_3_200 = 1.86e-05  mcrdlm5m1_cc_w_1_600_s_3_200 = 3.17e-11  mcrdlm5m1_cf_w_1_600_s_3_200 = 2.49e-11
+ mcrdlm5m1_ca_w_1_600_s_4_800 = 1.86e-05  mcrdlm5m1_cc_w_1_600_s_4_800 = 1.70e-11  mcrdlm5m1_cf_w_1_600_s_4_800 = 3.33e-11
+ mcrdlm5m1_ca_w_1_600_s_10_000 = 1.86e-05  mcrdlm5m1_cc_w_1_600_s_10_000 = 2.71e-12  mcrdlm5m1_cf_w_1_600_s_10_000 = 4.49e-11
+ mcrdlm5m1_ca_w_1_600_s_12_000 = 1.86e-05  mcrdlm5m1_cc_w_1_600_s_12_000 = 1.34e-12  mcrdlm5m1_cf_w_1_600_s_12_000 = 4.62e-11
+ mcrdlm5m1_ca_w_4_000_s_1_600 = 1.86e-05  mcrdlm5m1_cc_w_4_000_s_1_600 = 7.44e-11  mcrdlm5m1_cf_w_4_000_s_1_600 = 1.33e-11
+ mcrdlm5m1_ca_w_4_000_s_1_700 = 1.86e-05  mcrdlm5m1_cc_w_4_000_s_1_700 = 6.94e-11  mcrdlm5m1_cf_w_4_000_s_1_700 = 1.41e-11
+ mcrdlm5m1_ca_w_4_000_s_1_900 = 1.86e-05  mcrdlm5m1_cc_w_4_000_s_1_900 = 6.14e-11  mcrdlm5m1_cf_w_4_000_s_1_900 = 1.57e-11
+ mcrdlm5m1_ca_w_4_000_s_2_000 = 1.86e-05  mcrdlm5m1_cc_w_4_000_s_2_000 = 5.79e-11  mcrdlm5m1_cf_w_4_000_s_2_000 = 1.65e-11
+ mcrdlm5m1_ca_w_4_000_s_2_400 = 1.86e-05  mcrdlm5m1_cc_w_4_000_s_2_400 = 4.68e-11  mcrdlm5m1_cf_w_4_000_s_2_400 = 1.95e-11
+ mcrdlm5m1_ca_w_4_000_s_2_800 = 1.86e-05  mcrdlm5m1_cc_w_4_000_s_2_800 = 3.87e-11  mcrdlm5m1_cf_w_4_000_s_2_800 = 2.23e-11
+ mcrdlm5m1_ca_w_4_000_s_3_200 = 1.86e-05  mcrdlm5m1_cc_w_4_000_s_3_200 = 3.25e-11  mcrdlm5m1_cf_w_4_000_s_3_200 = 2.50e-11
+ mcrdlm5m1_ca_w_4_000_s_4_800 = 1.86e-05  mcrdlm5m1_cc_w_4_000_s_4_800 = 1.75e-11  mcrdlm5m1_cf_w_4_000_s_4_800 = 3.35e-11
+ mcrdlm5m1_ca_w_4_000_s_10_000 = 1.86e-05  mcrdlm5m1_cc_w_4_000_s_10_000 = 2.81e-12  mcrdlm5m1_cf_w_4_000_s_10_000 = 4.53e-11
+ mcrdlm5m1_ca_w_4_000_s_12_000 = 1.86e-05  mcrdlm5m1_cc_w_4_000_s_12_000 = 1.41e-12  mcrdlm5m1_cf_w_4_000_s_12_000 = 4.67e-11
+ mcrdlm5m2_ca_w_1_600_s_1_600 = 2.07e-05  mcrdlm5m2_cc_w_1_600_s_1_600 = 7.09e-11  mcrdlm5m2_cf_w_1_600_s_1_600 = 1.48e-11
+ mcrdlm5m2_ca_w_1_600_s_1_700 = 2.07e-05  mcrdlm5m2_cc_w_1_600_s_1_700 = 6.61e-11  mcrdlm5m2_cf_w_1_600_s_1_700 = 1.56e-11
+ mcrdlm5m2_ca_w_1_600_s_1_900 = 2.07e-05  mcrdlm5m2_cc_w_1_600_s_1_900 = 5.82e-11  mcrdlm5m2_cf_w_1_600_s_1_900 = 1.74e-11
+ mcrdlm5m2_ca_w_1_600_s_2_000 = 2.07e-05  mcrdlm5m2_cc_w_1_600_s_2_000 = 5.48e-11  mcrdlm5m2_cf_w_1_600_s_2_000 = 1.82e-11
+ mcrdlm5m2_ca_w_1_600_s_2_400 = 2.07e-05  mcrdlm5m2_cc_w_1_600_s_2_400 = 4.39e-11  mcrdlm5m2_cf_w_1_600_s_2_400 = 2.15e-11
+ mcrdlm5m2_ca_w_1_600_s_2_800 = 2.07e-05  mcrdlm5m2_cc_w_1_600_s_2_800 = 3.61e-11  mcrdlm5m2_cf_w_1_600_s_2_800 = 2.45e-11
+ mcrdlm5m2_ca_w_1_600_s_3_200 = 2.07e-05  mcrdlm5m2_cc_w_1_600_s_3_200 = 3.00e-11  mcrdlm5m2_cf_w_1_600_s_3_200 = 2.73e-11
+ mcrdlm5m2_ca_w_1_600_s_4_800 = 2.07e-05  mcrdlm5m2_cc_w_1_600_s_4_800 = 1.56e-11  mcrdlm5m2_cf_w_1_600_s_4_800 = 3.60e-11
+ mcrdlm5m2_ca_w_1_600_s_10_000 = 2.07e-05  mcrdlm5m2_cc_w_1_600_s_10_000 = 2.16e-12  mcrdlm5m2_cf_w_1_600_s_10_000 = 4.71e-11
+ mcrdlm5m2_ca_w_1_600_s_12_000 = 2.07e-05  mcrdlm5m2_cc_w_1_600_s_12_000 = 1.01e-12  mcrdlm5m2_cf_w_1_600_s_12_000 = 4.82e-11
+ mcrdlm5m2_ca_w_4_000_s_1_600 = 2.07e-05  mcrdlm5m2_cc_w_4_000_s_1_600 = 7.25e-11  mcrdlm5m2_cf_w_4_000_s_1_600 = 1.47e-11
+ mcrdlm5m2_ca_w_4_000_s_1_700 = 2.07e-05  mcrdlm5m2_cc_w_4_000_s_1_700 = 6.75e-11  mcrdlm5m2_cf_w_4_000_s_1_700 = 1.56e-11
+ mcrdlm5m2_ca_w_4_000_s_1_900 = 2.07e-05  mcrdlm5m2_cc_w_4_000_s_1_900 = 5.94e-11  mcrdlm5m2_cf_w_4_000_s_1_900 = 1.74e-11
+ mcrdlm5m2_ca_w_4_000_s_2_000 = 2.07e-05  mcrdlm5m2_cc_w_4_000_s_2_000 = 5.60e-11  mcrdlm5m2_cf_w_4_000_s_2_000 = 1.82e-11
+ mcrdlm5m2_ca_w_4_000_s_2_400 = 2.07e-05  mcrdlm5m2_cc_w_4_000_s_2_400 = 4.49e-11  mcrdlm5m2_cf_w_4_000_s_2_400 = 2.15e-11
+ mcrdlm5m2_ca_w_4_000_s_2_800 = 2.07e-05  mcrdlm5m2_cc_w_4_000_s_2_800 = 3.68e-11  mcrdlm5m2_cf_w_4_000_s_2_800 = 2.45e-11
+ mcrdlm5m2_ca_w_4_000_s_3_200 = 2.07e-05  mcrdlm5m2_cc_w_4_000_s_3_200 = 3.07e-11  mcrdlm5m2_cf_w_4_000_s_3_200 = 2.73e-11
+ mcrdlm5m2_ca_w_4_000_s_4_800 = 2.07e-05  mcrdlm5m2_cc_w_4_000_s_4_800 = 1.59e-11  mcrdlm5m2_cf_w_4_000_s_4_800 = 3.62e-11
+ mcrdlm5m2_ca_w_4_000_s_10_000 = 2.07e-05  mcrdlm5m2_cc_w_4_000_s_10_000 = 2.21e-12  mcrdlm5m2_cf_w_4_000_s_10_000 = 4.76e-11
+ mcrdlm5m2_ca_w_4_000_s_12_000 = 2.07e-05  mcrdlm5m2_cc_w_4_000_s_12_000 = 1.06e-12  mcrdlm5m2_cf_w_4_000_s_12_000 = 4.87e-11
+ mcrdlm5m3_ca_w_1_600_s_1_600 = 3.09e-05  mcrdlm5m3_cc_w_1_600_s_1_600 = 6.49e-11  mcrdlm5m3_cf_w_1_600_s_1_600 = 2.12e-11
+ mcrdlm5m3_ca_w_1_600_s_1_700 = 3.09e-05  mcrdlm5m3_cc_w_1_600_s_1_700 = 6.02e-11  mcrdlm5m3_cf_w_1_600_s_1_700 = 2.24e-11
+ mcrdlm5m3_ca_w_1_600_s_1_900 = 3.09e-05  mcrdlm5m3_cc_w_1_600_s_1_900 = 5.21e-11  mcrdlm5m3_cf_w_1_600_s_1_900 = 2.48e-11
+ mcrdlm5m3_ca_w_1_600_s_2_000 = 3.09e-05  mcrdlm5m3_cc_w_1_600_s_2_000 = 4.87e-11  mcrdlm5m3_cf_w_1_600_s_2_000 = 2.59e-11
+ mcrdlm5m3_ca_w_1_600_s_2_400 = 3.09e-05  mcrdlm5m3_cc_w_1_600_s_2_400 = 3.79e-11  mcrdlm5m3_cf_w_1_600_s_2_400 = 3.01e-11
+ mcrdlm5m3_ca_w_1_600_s_2_800 = 3.09e-05  mcrdlm5m3_cc_w_1_600_s_2_800 = 3.03e-11  mcrdlm5m3_cf_w_1_600_s_2_800 = 3.39e-11
+ mcrdlm5m3_ca_w_1_600_s_3_200 = 3.09e-05  mcrdlm5m3_cc_w_1_600_s_3_200 = 2.45e-11  mcrdlm5m3_cf_w_1_600_s_3_200 = 3.73e-11
+ mcrdlm5m3_ca_w_1_600_s_4_800 = 3.09e-05  mcrdlm5m3_cc_w_1_600_s_4_800 = 1.11e-11  mcrdlm5m3_cf_w_1_600_s_4_800 = 4.67e-11
+ mcrdlm5m3_ca_w_1_600_s_10_000 = 3.09e-05  mcrdlm5m3_cc_w_1_600_s_10_000 = 1.08e-12  mcrdlm5m3_cf_w_1_600_s_10_000 = 5.58e-11
+ mcrdlm5m3_ca_w_1_600_s_12_000 = 3.09e-05  mcrdlm5m3_cc_w_1_600_s_12_000 = 4.35e-13  mcrdlm5m3_cf_w_1_600_s_12_000 = 5.64e-11
+ mcrdlm5m3_ca_w_4_000_s_1_600 = 3.09e-05  mcrdlm5m3_cc_w_4_000_s_1_600 = 6.62e-11  mcrdlm5m3_cf_w_4_000_s_1_600 = 2.12e-11
+ mcrdlm5m3_ca_w_4_000_s_1_700 = 3.09e-05  mcrdlm5m3_cc_w_4_000_s_1_700 = 6.12e-11  mcrdlm5m3_cf_w_4_000_s_1_700 = 2.24e-11
+ mcrdlm5m3_ca_w_4_000_s_1_900 = 3.09e-05  mcrdlm5m3_cc_w_4_000_s_1_900 = 5.30e-11  mcrdlm5m3_cf_w_4_000_s_1_900 = 2.48e-11
+ mcrdlm5m3_ca_w_4_000_s_2_000 = 3.09e-05  mcrdlm5m3_cc_w_4_000_s_2_000 = 4.96e-11  mcrdlm5m3_cf_w_4_000_s_2_000 = 2.59e-11
+ mcrdlm5m3_ca_w_4_000_s_2_400 = 3.09e-05  mcrdlm5m3_cc_w_4_000_s_2_400 = 3.88e-11  mcrdlm5m3_cf_w_4_000_s_2_400 = 3.01e-11
+ mcrdlm5m3_ca_w_4_000_s_2_800 = 3.09e-05  mcrdlm5m3_cc_w_4_000_s_2_800 = 3.10e-11  mcrdlm5m3_cf_w_4_000_s_2_800 = 3.40e-11
+ mcrdlm5m3_ca_w_4_000_s_3_200 = 3.09e-05  mcrdlm5m3_cc_w_4_000_s_3_200 = 2.50e-11  mcrdlm5m3_cf_w_4_000_s_3_200 = 3.73e-11
+ mcrdlm5m3_ca_w_4_000_s_4_800 = 3.09e-05  mcrdlm5m3_cc_w_4_000_s_4_800 = 1.15e-11  mcrdlm5m3_cf_w_4_000_s_4_800 = 4.69e-11
+ mcrdlm5m3_ca_w_4_000_s_10_000 = 3.09e-05  mcrdlm5m3_cc_w_4_000_s_10_000 = 1.09e-12  mcrdlm5m3_cf_w_4_000_s_10_000 = 5.61e-11
+ mcrdlm5m3_ca_w_4_000_s_12_000 = 3.09e-05  mcrdlm5m3_cc_w_4_000_s_12_000 = 4.35e-13  mcrdlm5m3_cf_w_4_000_s_12_000 = 5.68e-11
+ mcrdlm5m4_ca_w_1_600_s_1_600 = 1.04e-04  mcrdlm5m4_cc_w_1_600_s_1_600 = 5.02e-11  mcrdlm5m4_cf_w_1_600_s_1_600 = 5.24e-11
+ mcrdlm5m4_ca_w_1_600_s_1_700 = 1.04e-04  mcrdlm5m4_cc_w_1_600_s_1_700 = 4.55e-11  mcrdlm5m4_cf_w_1_600_s_1_700 = 5.46e-11
+ mcrdlm5m4_ca_w_1_600_s_1_900 = 1.04e-04  mcrdlm5m4_cc_w_1_600_s_1_900 = 3.80e-11  mcrdlm5m4_cf_w_1_600_s_1_900 = 5.84e-11
+ mcrdlm5m4_ca_w_1_600_s_2_000 = 1.04e-04  mcrdlm5m4_cc_w_1_600_s_2_000 = 3.49e-11  mcrdlm5m4_cf_w_1_600_s_2_000 = 6.01e-11
+ mcrdlm5m4_ca_w_1_600_s_2_400 = 1.04e-04  mcrdlm5m4_cc_w_1_600_s_2_400 = 2.53e-11  mcrdlm5m4_cf_w_1_600_s_2_400 = 6.60e-11
+ mcrdlm5m4_ca_w_1_600_s_2_800 = 1.04e-04  mcrdlm5m4_cc_w_1_600_s_2_800 = 1.89e-11  mcrdlm5m4_cf_w_1_600_s_2_800 = 7.07e-11
+ mcrdlm5m4_ca_w_1_600_s_3_200 = 1.04e-04  mcrdlm5m4_cc_w_1_600_s_3_200 = 1.43e-11  mcrdlm5m4_cf_w_1_600_s_3_200 = 7.44e-11
+ mcrdlm5m4_ca_w_1_600_s_4_800 = 1.04e-04  mcrdlm5m4_cc_w_1_600_s_4_800 = 5.13e-12  mcrdlm5m4_cf_w_1_600_s_4_800 = 8.23e-11
+ mcrdlm5m4_ca_w_1_600_s_10_000 = 1.04e-04  mcrdlm5m4_cc_w_1_600_s_10_000 = 2.60e-13  mcrdlm5m4_cf_w_1_600_s_10_000 = 8.72e-11
+ mcrdlm5m4_ca_w_1_600_s_12_000 = 1.04e-04  mcrdlm5m4_cc_w_1_600_s_12_000 = 1.25e-13  mcrdlm5m4_cf_w_1_600_s_12_000 = 8.74e-11
+ mcrdlm5m4_ca_w_4_000_s_1_600 = 1.04e-04  mcrdlm5m4_cc_w_4_000_s_1_600 = 5.13e-11  mcrdlm5m4_cf_w_4_000_s_1_600 = 5.24e-11
+ mcrdlm5m4_ca_w_4_000_s_1_700 = 1.04e-04  mcrdlm5m4_cc_w_4_000_s_1_700 = 4.65e-11  mcrdlm5m4_cf_w_4_000_s_1_700 = 5.45e-11
+ mcrdlm5m4_ca_w_4_000_s_1_900 = 1.04e-04  mcrdlm5m4_cc_w_4_000_s_1_900 = 3.90e-11  mcrdlm5m4_cf_w_4_000_s_1_900 = 5.83e-11
+ mcrdlm5m4_ca_w_4_000_s_2_000 = 1.04e-04  mcrdlm5m4_cc_w_4_000_s_2_000 = 3.58e-11  mcrdlm5m4_cf_w_4_000_s_2_000 = 6.01e-11
+ mcrdlm5m4_ca_w_4_000_s_2_400 = 1.04e-04  mcrdlm5m4_cc_w_4_000_s_2_400 = 2.60e-11  mcrdlm5m4_cf_w_4_000_s_2_400 = 6.61e-11
+ mcrdlm5m4_ca_w_4_000_s_2_800 = 1.04e-04  mcrdlm5m4_cc_w_4_000_s_2_800 = 1.95e-11  mcrdlm5m4_cf_w_4_000_s_2_800 = 7.08e-11
+ mcrdlm5m4_ca_w_4_000_s_3_200 = 1.04e-04  mcrdlm5m4_cc_w_4_000_s_3_200 = 1.48e-11  mcrdlm5m4_cf_w_4_000_s_3_200 = 7.45e-11
+ mcrdlm5m4_ca_w_4_000_s_4_800 = 1.04e-04  mcrdlm5m4_cc_w_4_000_s_4_800 = 5.36e-12  mcrdlm5m4_cf_w_4_000_s_4_800 = 8.26e-11
+ mcrdlm5m4_ca_w_4_000_s_10_000 = 1.04e-04  mcrdlm5m4_cc_w_4_000_s_10_000 = 3.15e-13  mcrdlm5m4_cf_w_4_000_s_10_000 = 8.77e-11
+ mcrdlm5m4_ca_w_4_000_s_12_000 = 1.04e-04  mcrdlm5m4_cc_w_4_000_s_12_000 = 1.20e-13  mcrdlm5m4_cf_w_4_000_s_12_000 = 8.79e-11
+ cp1f = 1.36e-04  cp1fsw = 9.70e-11
+ cl1f = 4.51e-05  cl1fsw = 9.71e-11
+ cl1d = 6.56e-05  cl1dsw = 9.61e-11
+ cl1p1 = 1.40e-04  cl1p1sw = 9.46e-11
+ cm1f = 3.18e-05  cm1fsw = 1.24e-10
+ cm1d = 4.07e-05  cm1dsw = 1.24e-10
+ cm1p1 = 6.07e-05  cm1p1sw = 1.23e-10
+ cm1l1 = 1.63e-04  cm1l1sw = 1.18e-10
+ cm2f = 2.13e-05  cm2fsw = 1.25e-10
+ cm2d = 2.49e-05  cm2dsw = 1.24e-10
+ cm2p1 = 3.12e-05  cm2p1sw = 1.24e-10
+ cm2l1 = 4.60e-05  cm2l1sw = 1.23e-10
+ cm2m1 = 2.18e-04  cm2m1sw = 1.19e-10
+ cm3f = 1.49e-05  cm3fsw = 1.20e-10
+ cm3d = 1.67e-05  cm3dsw = 1.20e-10
+ cm3p1 = 1.92e-05  cm3p1sw = 1.20e-10
+ cm3l1 = 2.40e-05  cm3l1sw = 1.19e-10
+ cm3m1 = 4.08e-05  cm3m1sw = 1.18e-10
+ cm3m2 = 1.12e-04  cm3m2sw = 1.16e-10
+ cm4f = 9.99e-06  cm4fsw = 1.22e-10
+ cm4d = 1.07e-05  cm4dsw = 1.22e-10
+ cm4p1 = 1.17e-05  cm4p1sw = 1.22e-10
+ cm4l1 = 1.34e-05  cm4l1sw = 1.22e-10
+ cm4m1 = 1.73e-05  cm4m1sw = 1.21e-10
+ cm4m2 = 2.38e-05  cm4m2sw = 1.21e-10
+ cm4m3 = 1.42e-04  cm4m3sw = 1.18e-10
+ cm5f = 7.33e-06  cm5fsw = 9.03e-11
+ cm5d = 7.72e-06  cm5dsw = 9.01e-11
+ cm5p1 = 8.24e-06  cm5p1sw = 9.01e-11
+ cm5l1 = 8.99e-06  cm5l1sw = 9.00e-11
+ cm5m1 = 1.06e-05  cm5m1sw = 8.96e-11
+ cm5m2 = 1.27e-05  cm5m2sw = 8.94e-11
+ cm5m3 = 2.30e-05  cm5m3sw = 8.96e-11
+ cm5m4 = 9.63e-05  cm5m4sw = 1.06e-10
+ crdlf = 3.26e-06  crdlfsw = 7.06e-11
+ crdld = 3.34e-06  crdldsw = 7.05e-11
+ crdlp1 = 3.43e-06  crdlp1sw = 7.04e-11
+ crdll1 = 3.55e-06  crdll1sw = 7.03e-11
+ crdlm1 = 3.79e-06  crdlm1sw = 7.01e-11
+ crdlm2 = 4.02e-06  crdlm2sw = 6.99e-11
+ crdlm3 = 4.69e-06  crdlm3sw = 6.95e-11
+ crdlm4 = 5.55e-06  crdlm4sw = 6.92e-11
+ crdlm5 = 7.92e-06  crdlm5sw = 6.95e-11
+ cl1p1f = 2.76e-04  cl1p1fsw = 9.25e-11
+ cm1p1f = 1.97e-04  cm1p1fsw = 9.41e-11
+ cm2p1f = 1.67e-04  cm2p1fsw = 9.55e-11
+ cm3p1f = 1.55e-04  cm3p1fsw = 9.62e-11
+ cm4p1f = 1.48e-04  cm4p1fsw = 9.65e-11
+ cm5p1f = 1.44e-04  cm5p1fsw = 9.67e-11
+ crdlp1f = 1.39e-04  crdlp1fsw = 9.69e-11
+ cm1l1f = 2.08e-04  cm1l1fsw = 9.10e-11
+ cm1l1d = 2.29e-04  cm1l1dsw = 9.01e-11
+ cm1l1p1 = 3.04e-04  cm1l1p1sw = 8.85e-11
+ cm2l1f = 9.12e-05  cm2l1fsw = 9.38e-11
+ cm2l1d = 1.12e-04  cm2l1dsw = 9.28e-11
+ cm2l1p1 = 1.86e-04  cm2l1p1sw = 9.17e-11
+ cm3l1f = 6.92e-05  cm3l1fsw = 9.53e-11
+ cm3l1d = 8.97e-05  cm3l1dsw = 9.43e-11
+ cm3l1p1 = 1.64e-04  cm3l1p1sw = 9.31e-11
+ cm4l1f = 5.85e-05  cm4l1fsw = 9.60e-11
+ cm4l1d = 7.90e-05  cm4l1dsw = 9.51e-11
+ cm4l1p1 = 1.53e-04  cm4l1p1sw = 9.38e-11
+ cm5l1f = 5.41e-05  cm5l1fsw = 9.63e-11
+ cm5l1d = 7.46e-05  cm5l1dsw = 9.54e-11
+ cm5l1p1 = 1.49e-04  cm5l1p1sw = 9.41e-11
+ crdll1f = 4.87e-05  crdll1fsw = 9.66e-11
+ crdll1d = 6.92e-05  crdll1dsw = 9.59e-11
+ crdll1p1 = 1.44e-04  crdll1p1sw = 9.44e-11
+ cm2m1f = 2.50e-04  cm2m1fsw = 1.16e-10
+ cm2m1d = 2.59e-04  cm2m1dsw = 1.16e-10
+ cm2m1p1 = 2.79e-04  cm2m1p1sw = 1.16e-10
+ cm2m1l1 = 3.81e-04  cm2m1l1sw = 1.12e-10
+ cm3m1f = 7.26e-05  cm3m1fsw = 1.21e-10
+ cm3m1d = 8.16e-05  cm3m1dsw = 1.20e-10
+ cm3m1p1 = 1.02e-04  cm3m1p1sw = 1.18e-10
+ cm3m1l1 = 2.04e-04  cm3m1l1sw = 1.17e-10
+ cm4m1f = 4.91e-05  cm4m1fsw = 1.23e-10
+ cm4m1d = 5.81e-05  cm4m1dsw = 1.21e-10
+ cm4m1p1 = 7.81e-05  cm4m1p1sw = 1.20e-10
+ cm4m1l1 = 1.80e-04  cm4m1l1sw = 1.18e-10
+ cm5m1f = 4.24e-05  cm5m1fsw = 1.23e-10
+ cm5m1d = 5.14e-05  cm5m1dsw = 1.21e-10
+ cm5m1p1 = 7.14e-05  cm5m1p1sw = 1.20e-10
+ cm5m1l1 = 1.73e-04  cm5m1l1sw = 1.19e-10
+ crdlm1f = 3.56e-05  crdlm1fsw = 1.24e-10
+ crdlm1d = 4.45e-05  crdlm1dsw = 1.21e-10
+ crdlm1p1 = 6.45e-05  crdlm1p1sw = 1.20e-10
+ crdlm1l1 = 1.67e-04  crdlm1l1sw = 1.18e-10
+ cm3m2f = 1.34e-04  cm3m2fsw = 1.18e-10
+ cm3m2d = 1.37e-04  cm3m2dsw = 1.18e-10
+ cm3m2p1 = 1.44e-04  cm3m2p1sw = 1.17e-10
+ cm3m2l1 = 1.58e-04  cm3m2l1sw = 1.17e-10
+ cm3m2m1 = 3.31e-04  cm3m2m1sw = 1.13e-10
+ cm4m2f = 4.50e-05  cm4m2fsw = 1.23e-10
+ cm4m2d = 4.87e-05  cm4m2dsw = 1.22e-10
+ cm4m2p1 = 5.50e-05  cm4m2p1sw = 1.21e-10
+ cm4m2l1 = 6.98e-05  cm4m2l1sw = 1.20e-10
+ cm4m2m1 = 2.42e-04  cm4m2m1sw = 1.18e-10
+ cm5m2f = 3.40e-05  cm5m2fsw = 1.23e-10
+ cm5m2d = 3.77e-05  cm5m2dsw = 1.23e-10
+ cm5m2p1 = 4.39e-05  cm5m2p1sw = 1.21e-10
+ cm5m2l1 = 5.87e-05  cm5m2l1sw = 1.20e-10
+ cm5m2m1 = 2.31e-04  cm5m2m1sw = 1.18e-10
+ crdlm2f = 2.53e-05  crdlm2fsw = 1.24e-10
+ crdlm2d = 2.89e-05  crdlm2dsw = 1.23e-10
+ crdlm2p1 = 3.52e-05  crdlm2p1sw = 1.21e-10
+ crdlm2l1 = 5.00e-05  crdlm2l1sw = 1.21e-10
+ crdlm2m1 = 2.22e-04  crdlm2m1sw = 1.19e-10
+ cm4m3f = 1.57e-04  cm4m3fsw = 1.14e-10
+ cm4m3d = 1.59e-04  cm4m3dsw = 1.14e-10
+ cm4m3p1 = 1.61e-04  cm4m3p1sw = 1.14e-10
+ cm4m3l1 = 1.66e-04  cm4m3l1sw = 1.13e-10
+ cm4m3m1 = 1.83e-04  cm4m3m1sw = 1.12e-10
+ cm4m3m2 = 2.54e-04  cm4m3m2sw = 1.10e-10
+ cm5m3f = 3.79e-05  cm5m3fsw = 1.18e-10
+ cm5m3d = 3.96e-05  cm5m3dsw = 1.18e-10
+ cm5m3p1 = 4.22e-05  cm5m3p1sw = 1.17e-10
+ cm5m3l1 = 4.70e-05  cm5m3l1sw = 1.17e-10
+ cm5m3m1 = 6.38e-05  cm5m3m1sw = 1.15e-10
+ cm5m3m2 = 1.35e-04  cm5m3m2sw = 1.14e-10
+ crdlm3f = 1.96e-05  crdlm3fsw = 1.20e-10
+ crdlm3d = 2.13e-05  crdlm3dsw = 1.20e-10
+ crdlm3p1 = 2.39e-05  crdlm3p1sw = 1.19e-10
+ crdlm3l1 = 2.87e-05  crdlm3l1sw = 1.19e-10
+ crdlm3m1 = 4.55e-05  crdlm3m1sw = 1.18e-10
+ crdlm3m2 = 1.17e-04  crdlm3m2sw = 1.16e-10
+ cm5m4f = 1.06e-04  cm5m4fsw = 1.14e-10
+ cm5m4d = 1.07e-04  cm5m4dsw = 1.14e-10
+ cm5m4p1 = 1.08e-04  cm5m4p1sw = 1.14e-10
+ cm5m4l1 = 1.10e-04  cm5m4l1sw = 1.14e-10
+ cm5m4m1 = 1.14e-04  cm5m4m1sw = 1.14e-10
+ cm5m4m2 = 1.20e-04  cm5m4m2sw = 1.13e-10
+ cm5m4m3 = 2.38e-04  cm5m4m3sw = 1.11e-10
+ crdlm4f = 1.55e-05  crdlm4fsw = 1.22e-10
+ crdlm4d = 1.63e-05  crdlm4dsw = 1.22e-10
+ crdlm4p1 = 1.73e-05  crdlm4p1sw = 1.21e-10
+ crdlm4l1 = 1.89e-05  crdlm4l1sw = 1.21e-10
+ crdlm4m1 = 2.29e-05  crdlm4m1sw = 1.21e-10
+ crdlm4m2 = 2.93e-05  crdlm4m2sw = 1.20e-10
+ crdlm4m3 = 1.47e-04  crdlm4m3sw = 1.18e-10
+ crdlm5f = 1.53e-05  crdlm5fsw = 8.66e-11
+ crdlm5d = 1.57e-05  crdlm5dsw = 8.65e-11
+ crdlm5p1 = 1.62e-05  crdlm5p1sw = 8.63e-11
+ crdlm5l1 = 1.69e-05  crdlm5l1sw = 8.63e-11
+ crdlm5m1 = 1.86e-05  crdlm5m1sw = 8.60e-11
+ crdlm5m2 = 2.07e-05  crdlm5m2sw = 8.57e-11
+ crdlm5m3 = 3.09e-05  crdlm5m3sw = 8.61e-11
+ crdlm5m4 = 1.04e-04  crdlm5m4sw = 1.03e-10
