* SKY130 Spice File.
