* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.

* SKY130 Spice File.
* Number of bins: 52
.param
+ sky130_fd_pr__pfet_01v8__toxe_mult = 0.948
+ sky130_fd_pr__pfet_01v8__rshp_mult = 1.0
+ sky130_fd_pr__pfet_01v8__overlap_mult = 0.95436
+ sky130_fd_pr__pfet_01v8__ajunction_mult = 0.90161
+ sky130_fd_pr__pfet_01v8__pjunction_mult = 0.90587
+ sky130_fd_pr__pfet_01v8__lint_diff = 1.7325e-8
+ sky130_fd_pr__pfet_01v8__wint_diff = -3.2175e-8
+ sky130_fd_pr__pfet_01v8__dlc_diff = 1.7325e-8
+ sky130_fd_pr__pfet_01v8__dwc_diff = -3.2175e-8
*
* sky130_fd_pr__pfet_01v8, Bin 000, W = 1.26, L = 0.15
* -----------------------------------
+ sky130_fd_pr__pfet_01v8__agidl_diff_0 = 0.0
+ sky130_fd_pr__pfet_01v8__nfactor_diff_0 = 2.7052
+ sky130_fd_pr__pfet_01v8__vsat_diff_0 = -13041.0
+ sky130_fd_pr__pfet_01v8__a0_diff_0 = 0.0
+ sky130_fd_pr__pfet_01v8__pdits_diff_0 = 0.0
+ sky130_fd_pr__pfet_01v8__b0_diff_0 = 0.0
+ sky130_fd_pr__pfet_01v8__pclm_diff_0 = 0.0
+ sky130_fd_pr__pfet_01v8__kt1_diff_0 = 0.0
+ sky130_fd_pr__pfet_01v8__eta0_diff_0 = 0.0
+ sky130_fd_pr__pfet_01v8__ua_diff_0 = -2.3326e-12
+ sky130_fd_pr__pfet_01v8__keta_diff_0 = 0.0
+ sky130_fd_pr__pfet_01v8__rdsw_diff_0 = 0.0
+ sky130_fd_pr__pfet_01v8__k2_diff_0 = 0.0045512
+ sky130_fd_pr__pfet_01v8__vth0_diff_0 = -0.054958
+ sky130_fd_pr__pfet_01v8__pditsd_diff_0 = 0.0
+ sky130_fd_pr__pfet_01v8__u0_diff_0 = 0.00064676
+ sky130_fd_pr__pfet_01v8__b1_diff_0 = 0.0
+ sky130_fd_pr__pfet_01v8__cgidl_diff_0 = 0.0
+ sky130_fd_pr__pfet_01v8__tvoff_diff_0 = 0.0
+ sky130_fd_pr__pfet_01v8__voff_diff_0 = -0.23485
+ sky130_fd_pr__pfet_01v8__ags_diff_0 = 0.0
+ sky130_fd_pr__pfet_01v8__bgidl_diff_0 = 0.0
+ sky130_fd_pr__pfet_01v8__ub_diff_0 = 4.1498e-19
*
* sky130_fd_pr__pfet_01v8, Bin 001, W = 1.68, L = 0.15
* -----------------------------------
+ sky130_fd_pr__pfet_01v8__bgidl_diff_1 = 0.0
+ sky130_fd_pr__pfet_01v8__ub_diff_1 = 3.0525e-19
+ sky130_fd_pr__pfet_01v8__agidl_diff_1 = 0.0
+ sky130_fd_pr__pfet_01v8__nfactor_diff_1 = 2.678
+ sky130_fd_pr__pfet_01v8__vsat_diff_1 = -16028.0
+ sky130_fd_pr__pfet_01v8__a0_diff_1 = 0.0
+ sky130_fd_pr__pfet_01v8__pdits_diff_1 = 0.0
+ sky130_fd_pr__pfet_01v8__b0_diff_1 = 0.0
+ sky130_fd_pr__pfet_01v8__pclm_diff_1 = 0.0
+ sky130_fd_pr__pfet_01v8__kt1_diff_1 = 0.0
+ sky130_fd_pr__pfet_01v8__eta0_diff_1 = 0.0
+ sky130_fd_pr__pfet_01v8__ua_diff_1 = -3.8211e-11
+ sky130_fd_pr__pfet_01v8__keta_diff_1 = 0.0
+ sky130_fd_pr__pfet_01v8__rdsw_diff_1 = 0.0
+ sky130_fd_pr__pfet_01v8__k2_diff_1 = 4.4689e-5
+ sky130_fd_pr__pfet_01v8__vth0_diff_1 = -0.1267
+ sky130_fd_pr__pfet_01v8__pditsd_diff_1 = 0.0
+ sky130_fd_pr__pfet_01v8__u0_diff_1 = 0.0003497
+ sky130_fd_pr__pfet_01v8__b1_diff_1 = 0.0
+ sky130_fd_pr__pfet_01v8__cgidl_diff_1 = 0.0
+ sky130_fd_pr__pfet_01v8__tvoff_diff_1 = 0.0
+ sky130_fd_pr__pfet_01v8__voff_diff_1 = -0.20996
+ sky130_fd_pr__pfet_01v8__ags_diff_1 = 0.0
*
* sky130_fd_pr__pfet_01v8, Bin 002, W = 1.0, L = 1.0
* ---------------------------------
+ sky130_fd_pr__pfet_01v8__cgidl_diff_2 = 0.0
+ sky130_fd_pr__pfet_01v8__tvoff_diff_2 = 0.0
+ sky130_fd_pr__pfet_01v8__voff_diff_2 = -0.097678
+ sky130_fd_pr__pfet_01v8__ags_diff_2 = -0.002113
+ sky130_fd_pr__pfet_01v8__bgidl_diff_2 = 0.0
+ sky130_fd_pr__pfet_01v8__ub_diff_2 = 5.467e-19
+ sky130_fd_pr__pfet_01v8__agidl_diff_2 = 0.0
+ sky130_fd_pr__pfet_01v8__nfactor_diff_2 = 0.15089
+ sky130_fd_pr__pfet_01v8__vsat_diff_2 = 0.0
+ sky130_fd_pr__pfet_01v8__a0_diff_2 = 0.0021271
+ sky130_fd_pr__pfet_01v8__pdits_diff_2 = 0.0
+ sky130_fd_pr__pfet_01v8__b0_diff_2 = 0.0
+ sky130_fd_pr__pfet_01v8__pclm_diff_2 = 0.0
+ sky130_fd_pr__pfet_01v8__kt1_diff_2 = 0.0
+ sky130_fd_pr__pfet_01v8__eta0_diff_2 = 0.0
+ sky130_fd_pr__pfet_01v8__ua_diff_2 = 3.5075e-12
+ sky130_fd_pr__pfet_01v8__keta_diff_2 = 0.0
+ sky130_fd_pr__pfet_01v8__rdsw_diff_2 = 0.0
+ sky130_fd_pr__pfet_01v8__k2_diff_2 = -0.0075788
+ sky130_fd_pr__pfet_01v8__vth0_diff_2 = 0.016199
+ sky130_fd_pr__pfet_01v8__pditsd_diff_2 = 0.0
+ sky130_fd_pr__pfet_01v8__u0_diff_2 = 0.0023435
+ sky130_fd_pr__pfet_01v8__b1_diff_2 = 0.0
*
* sky130_fd_pr__pfet_01v8, Bin 003, W = 1.0, L = 2.0
* ---------------------------------
+ sky130_fd_pr__pfet_01v8__b1_diff_3 = 0.0
+ sky130_fd_pr__pfet_01v8__cgidl_diff_3 = 0.0
+ sky130_fd_pr__pfet_01v8__tvoff_diff_3 = 0.0
+ sky130_fd_pr__pfet_01v8__voff_diff_3 = -0.10546
+ sky130_fd_pr__pfet_01v8__ags_diff_3 = -0.0036028
+ sky130_fd_pr__pfet_01v8__bgidl_diff_3 = 0.0
+ sky130_fd_pr__pfet_01v8__ub_diff_3 = 6.3506e-19
+ sky130_fd_pr__pfet_01v8__nfactor_diff_3 = 0.18478
+ sky130_fd_pr__pfet_01v8__vsat_diff_3 = 0.0
+ sky130_fd_pr__pfet_01v8__agidl_diff_3 = 0.0
+ sky130_fd_pr__pfet_01v8__a0_diff_3 = 0.0040252
+ sky130_fd_pr__pfet_01v8__pdits_diff_3 = 0.0
+ sky130_fd_pr__pfet_01v8__b0_diff_3 = 0.0
+ sky130_fd_pr__pfet_01v8__pclm_diff_3 = 0.0
+ sky130_fd_pr__pfet_01v8__kt1_diff_3 = 0.0
+ sky130_fd_pr__pfet_01v8__eta0_diff_3 = 0.0
+ sky130_fd_pr__pfet_01v8__ua_diff_3 = -2.4052e-12
+ sky130_fd_pr__pfet_01v8__keta_diff_3 = 0.0
+ sky130_fd_pr__pfet_01v8__rdsw_diff_3 = 0.0
+ sky130_fd_pr__pfet_01v8__k2_diff_3 = -0.012185
+ sky130_fd_pr__pfet_01v8__vth0_diff_3 = 0.021481
+ sky130_fd_pr__pfet_01v8__pditsd_diff_3 = 0.0
+ sky130_fd_pr__pfet_01v8__u0_diff_3 = 0.0028621
*
* sky130_fd_pr__pfet_01v8, Bin 004, W = 1.0, L = 4.0
* ---------------------------------
+ sky130_fd_pr__pfet_01v8__pditsd_diff_4 = 0.0
+ sky130_fd_pr__pfet_01v8__u0_diff_4 = 0.0029153
+ sky130_fd_pr__pfet_01v8__vth0_diff_4 = 0.0066881
+ sky130_fd_pr__pfet_01v8__b1_diff_4 = 0.0
+ sky130_fd_pr__pfet_01v8__cgidl_diff_4 = 0.0
+ sky130_fd_pr__pfet_01v8__tvoff_diff_4 = 0.0
+ sky130_fd_pr__pfet_01v8__voff_diff_4 = -0.10599
+ sky130_fd_pr__pfet_01v8__ags_diff_4 = 0.0051938
+ sky130_fd_pr__pfet_01v8__ub_diff_4 = 6.1783e-19
+ sky130_fd_pr__pfet_01v8__bgidl_diff_4 = 0.0
+ sky130_fd_pr__pfet_01v8__nfactor_diff_4 = 0.18255
+ sky130_fd_pr__pfet_01v8__vsat_diff_4 = 0.0
+ sky130_fd_pr__pfet_01v8__agidl_diff_4 = 0.0
+ sky130_fd_pr__pfet_01v8__a0_diff_4 = -0.0046292
+ sky130_fd_pr__pfet_01v8__pdits_diff_4 = 0.0
+ sky130_fd_pr__pfet_01v8__b0_diff_4 = 0.0
+ sky130_fd_pr__pfet_01v8__pclm_diff_4 = 0.0
+ sky130_fd_pr__pfet_01v8__kt1_diff_4 = 0.0
+ sky130_fd_pr__pfet_01v8__eta0_diff_4 = 0.0
+ sky130_fd_pr__pfet_01v8__ua_diff_4 = 3.5061e-13
+ sky130_fd_pr__pfet_01v8__keta_diff_4 = 0.0
+ sky130_fd_pr__pfet_01v8__rdsw_diff_4 = 0.0
+ sky130_fd_pr__pfet_01v8__k2_diff_4 = -0.013265
*
* sky130_fd_pr__pfet_01v8, Bin 005, W = 1.0, L = 8.0
* ---------------------------------
+ sky130_fd_pr__pfet_01v8__keta_diff_5 = 0.0
+ sky130_fd_pr__pfet_01v8__k2_diff_5 = -0.015073
+ sky130_fd_pr__pfet_01v8__pditsd_diff_5 = 0.0
+ sky130_fd_pr__pfet_01v8__u0_diff_5 = 0.0024177
+ sky130_fd_pr__pfet_01v8__vth0_diff_5 = -0.0092847
+ sky130_fd_pr__pfet_01v8__b1_diff_5 = 0.0
+ sky130_fd_pr__pfet_01v8__voff_diff_5 = -0.12061
+ sky130_fd_pr__pfet_01v8__cgidl_diff_5 = 0.0
+ sky130_fd_pr__pfet_01v8__tvoff_diff_5 = 0.0
+ sky130_fd_pr__pfet_01v8__ags_diff_5 = 0.049422
+ sky130_fd_pr__pfet_01v8__ub_diff_5 = 5.1769e-19
+ sky130_fd_pr__pfet_01v8__bgidl_diff_5 = 0.0
+ sky130_fd_pr__pfet_01v8__nfactor_diff_5 = 0.29986
+ sky130_fd_pr__pfet_01v8__vsat_diff_5 = 0.0
+ sky130_fd_pr__pfet_01v8__agidl_diff_5 = 0.0
+ sky130_fd_pr__pfet_01v8__a0_diff_5 = -0.045455
+ sky130_fd_pr__pfet_01v8__pdits_diff_5 = 0.0
+ sky130_fd_pr__pfet_01v8__b0_diff_5 = 0.0
+ sky130_fd_pr__pfet_01v8__pclm_diff_5 = 0.0
+ sky130_fd_pr__pfet_01v8__kt1_diff_5 = 0.0
+ sky130_fd_pr__pfet_01v8__eta0_diff_5 = 0.0
+ sky130_fd_pr__pfet_01v8__ua_diff_5 = -6.2498e-12
+ sky130_fd_pr__pfet_01v8__rdsw_diff_5 = 0.0
*
* sky130_fd_pr__pfet_01v8, Bin 006, W = 1.0, L = 0.15
* ----------------------------------
+ sky130_fd_pr__pfet_01v8__rdsw_diff_6 = 0.0
+ sky130_fd_pr__pfet_01v8__keta_diff_6 = 0.0
+ sky130_fd_pr__pfet_01v8__k2_diff_6 = 0.025127
+ sky130_fd_pr__pfet_01v8__pditsd_diff_6 = 0.0
+ sky130_fd_pr__pfet_01v8__u0_diff_6 = -0.00051028
+ sky130_fd_pr__pfet_01v8__vth0_diff_6 = -0.10272
+ sky130_fd_pr__pfet_01v8__b1_diff_6 = 0.0
+ sky130_fd_pr__pfet_01v8__voff_diff_6 = -0.16209
+ sky130_fd_pr__pfet_01v8__cgidl_diff_6 = 0.0
+ sky130_fd_pr__pfet_01v8__tvoff_diff_6 = 0.0
+ sky130_fd_pr__pfet_01v8__ags_diff_6 = 0.0
+ sky130_fd_pr__pfet_01v8__ub_diff_6 = 7.825e-19
+ sky130_fd_pr__pfet_01v8__bgidl_diff_6 = 0.0
+ sky130_fd_pr__pfet_01v8__nfactor_diff_6 = 2.176
+ sky130_fd_pr__pfet_01v8__vsat_diff_6 = -21227.0
+ sky130_fd_pr__pfet_01v8__agidl_diff_6 = 0.0
+ sky130_fd_pr__pfet_01v8__a0_diff_6 = 0.0
+ sky130_fd_pr__pfet_01v8__pdits_diff_6 = 0.0
+ sky130_fd_pr__pfet_01v8__b0_diff_6 = 0.0
+ sky130_fd_pr__pfet_01v8__pclm_diff_6 = 0.0
+ sky130_fd_pr__pfet_01v8__kt1_diff_6 = 0.0
+ sky130_fd_pr__pfet_01v8__eta0_diff_6 = 0.0
+ sky130_fd_pr__pfet_01v8__ua_diff_6 = -5.0e-10
*
* sky130_fd_pr__pfet_01v8, Bin 007, W = 1.0, L = 0.18
* ----------------------------------
+ sky130_fd_pr__pfet_01v8__kt1_diff_7 = 0.0
+ sky130_fd_pr__pfet_01v8__eta0_diff_7 = 0.0
+ sky130_fd_pr__pfet_01v8__ua_diff_7 = 1.2857e-10
+ sky130_fd_pr__pfet_01v8__rdsw_diff_7 = 0.0
+ sky130_fd_pr__pfet_01v8__keta_diff_7 = 0.0
+ sky130_fd_pr__pfet_01v8__k2_diff_7 = -0.00076543
+ sky130_fd_pr__pfet_01v8__pditsd_diff_7 = 0.0
+ sky130_fd_pr__pfet_01v8__u0_diff_7 = 0.00073453
+ sky130_fd_pr__pfet_01v8__vth0_diff_7 = -0.086522
+ sky130_fd_pr__pfet_01v8__b1_diff_7 = 0.0
+ sky130_fd_pr__pfet_01v8__voff_diff_7 = -0.26215
+ sky130_fd_pr__pfet_01v8__cgidl_diff_7 = 0.0
+ sky130_fd_pr__pfet_01v8__tvoff_diff_7 = 0.0
+ sky130_fd_pr__pfet_01v8__ags_diff_7 = 0.0
+ sky130_fd_pr__pfet_01v8__ub_diff_7 = 2.2283e-19
+ sky130_fd_pr__pfet_01v8__bgidl_diff_7 = 0.0
+ sky130_fd_pr__pfet_01v8__nfactor_diff_7 = 1.9904
+ sky130_fd_pr__pfet_01v8__vsat_diff_7 = -20000.0
+ sky130_fd_pr__pfet_01v8__agidl_diff_7 = 0.0
+ sky130_fd_pr__pfet_01v8__a0_diff_7 = 0.0
+ sky130_fd_pr__pfet_01v8__pdits_diff_7 = 0.0
+ sky130_fd_pr__pfet_01v8__b0_diff_7 = 0.0
+ sky130_fd_pr__pfet_01v8__pclm_diff_7 = 0.0
*
* sky130_fd_pr__pfet_01v8, Bin 008, W = 1.0, L = 0.25
* ----------------------------------
+ sky130_fd_pr__pfet_01v8__pclm_diff_8 = 0.0
+ sky130_fd_pr__pfet_01v8__kt1_diff_8 = 0.0
+ sky130_fd_pr__pfet_01v8__eta0_diff_8 = 0.0
+ sky130_fd_pr__pfet_01v8__ua_diff_8 = 2.7416e-11
+ sky130_fd_pr__pfet_01v8__rdsw_diff_8 = 0.0
+ sky130_fd_pr__pfet_01v8__keta_diff_8 = 0.0
+ sky130_fd_pr__pfet_01v8__k2_diff_8 = -0.0021971
+ sky130_fd_pr__pfet_01v8__pditsd_diff_8 = 0.0
+ sky130_fd_pr__pfet_01v8__u0_diff_8 = 4.347e-5
+ sky130_fd_pr__pfet_01v8__vth0_diff_8 = 0.028852
+ sky130_fd_pr__pfet_01v8__b1_diff_8 = 0.0
+ sky130_fd_pr__pfet_01v8__voff_diff_8 = -0.20736
+ sky130_fd_pr__pfet_01v8__cgidl_diff_8 = 0.0
+ sky130_fd_pr__pfet_01v8__tvoff_diff_8 = 0.0
+ sky130_fd_pr__pfet_01v8__ags_diff_8 = 0.0
+ sky130_fd_pr__pfet_01v8__ub_diff_8 = 2.9171e-19
+ sky130_fd_pr__pfet_01v8__bgidl_diff_8 = 0.0
+ sky130_fd_pr__pfet_01v8__nfactor_diff_8 = 1.1224
+ sky130_fd_pr__pfet_01v8__vsat_diff_8 = -11653.0
+ sky130_fd_pr__pfet_01v8__agidl_diff_8 = 0.0
+ sky130_fd_pr__pfet_01v8__a0_diff_8 = 0.0
+ sky130_fd_pr__pfet_01v8__pdits_diff_8 = 0.0
+ sky130_fd_pr__pfet_01v8__b0_diff_8 = 0.0
*
* sky130_fd_pr__pfet_01v8, Bin 009, W = 1.0, L = 0.5
* ---------------------------------
+ sky130_fd_pr__pfet_01v8__pdits_diff_9 = 0.0
+ sky130_fd_pr__pfet_01v8__b0_diff_9 = 0.0
+ sky130_fd_pr__pfet_01v8__pclm_diff_9 = 0.0
+ sky130_fd_pr__pfet_01v8__kt1_diff_9 = 0.0
+ sky130_fd_pr__pfet_01v8__eta0_diff_9 = 0.0
+ sky130_fd_pr__pfet_01v8__ua_diff_9 = 1.0972e-12
+ sky130_fd_pr__pfet_01v8__rdsw_diff_9 = 0.0
+ sky130_fd_pr__pfet_01v8__keta_diff_9 = 0.0
+ sky130_fd_pr__pfet_01v8__k2_diff_9 = -0.0087514
+ sky130_fd_pr__pfet_01v8__pditsd_diff_9 = 0.0
+ sky130_fd_pr__pfet_01v8__u0_diff_9 = 0.0011707
+ sky130_fd_pr__pfet_01v8__vth0_diff_9 = 0.044728
+ sky130_fd_pr__pfet_01v8__b1_diff_9 = 0.0
+ sky130_fd_pr__pfet_01v8__voff_diff_9 = -0.11579
+ sky130_fd_pr__pfet_01v8__cgidl_diff_9 = 0.0
+ sky130_fd_pr__pfet_01v8__tvoff_diff_9 = 0.0
+ sky130_fd_pr__pfet_01v8__ags_diff_9 = 0.0
+ sky130_fd_pr__pfet_01v8__ub_diff_9 = 4.4605e-19
+ sky130_fd_pr__pfet_01v8__bgidl_diff_9 = 0.0
+ sky130_fd_pr__pfet_01v8__nfactor_diff_9 = 0.27815
+ sky130_fd_pr__pfet_01v8__vsat_diff_9 = -3032.7
+ sky130_fd_pr__pfet_01v8__agidl_diff_9 = 0.0
+ sky130_fd_pr__pfet_01v8__a0_diff_9 = 0.0
*
* sky130_fd_pr__pfet_01v8, Bin 010, W = 2.0, L = 0.15
* ----------------------------------
+ sky130_fd_pr__pfet_01v8__pditsd_diff_10 = 0.0
+ sky130_fd_pr__pfet_01v8__eta0_diff_10 = 0.0
+ sky130_fd_pr__pfet_01v8__vsat_diff_10 = -20000.0
+ sky130_fd_pr__pfet_01v8__u0_diff_10 = -0.00070492
+ sky130_fd_pr__pfet_01v8__vth0_diff_10 = -0.086385
+ sky130_fd_pr__pfet_01v8__cgidl_diff_10 = 0.0
+ sky130_fd_pr__pfet_01v8__keta_diff_10 = 0.0
+ sky130_fd_pr__pfet_01v8__rdsw_diff_10 = 0.0
+ sky130_fd_pr__pfet_01v8__kt1_diff_10 = 0.0
+ sky130_fd_pr__pfet_01v8__pclm_diff_10 = 0.0
+ sky130_fd_pr__pfet_01v8__b0_diff_10 = 0.0
+ sky130_fd_pr__pfet_01v8__b1_diff_10 = 0.0
+ sky130_fd_pr__pfet_01v8__agidl_diff_10 = 0.0
+ sky130_fd_pr__pfet_01v8__ua_diff_10 = -2.9668e-10
+ sky130_fd_pr__pfet_01v8__bgidl_diff_10 = 0.0
+ sky130_fd_pr__pfet_01v8__nfactor_diff_10 = 1.2074
+ sky130_fd_pr__pfet_01v8__ub_diff_10 = 3.3082e-19
+ sky130_fd_pr__pfet_01v8__pdits_diff_10 = 0.0
+ sky130_fd_pr__pfet_01v8__tvoff_diff_10 = 0.0
+ sky130_fd_pr__pfet_01v8__ags_diff_10 = 0.0
+ sky130_fd_pr__pfet_01v8__k2_diff_10 = 0.039771
+ sky130_fd_pr__pfet_01v8__voff_diff_10 = -0.10113
+ sky130_fd_pr__pfet_01v8__a0_diff_10 = 0.0
*
* sky130_fd_pr__pfet_01v8, Bin 011, W = 3.0, L = 1.0
* ---------------------------------
+ sky130_fd_pr__pfet_01v8__voff_diff_11 = -0.11001
+ sky130_fd_pr__pfet_01v8__a0_diff_11 = -0.079538
+ sky130_fd_pr__pfet_01v8__pditsd_diff_11 = 0.0
+ sky130_fd_pr__pfet_01v8__eta0_diff_11 = 0.0
+ sky130_fd_pr__pfet_01v8__vsat_diff_11 = 27194.0
+ sky130_fd_pr__pfet_01v8__u0_diff_11 = 0.0018193
+ sky130_fd_pr__pfet_01v8__vth0_diff_11 = 0.0035882
+ sky130_fd_pr__pfet_01v8__cgidl_diff_11 = 0.0
+ sky130_fd_pr__pfet_01v8__keta_diff_11 = 0.0
+ sky130_fd_pr__pfet_01v8__rdsw_diff_11 = 0.0
+ sky130_fd_pr__pfet_01v8__kt1_diff_11 = 0.0
+ sky130_fd_pr__pfet_01v8__pclm_diff_11 = 0.0
+ sky130_fd_pr__pfet_01v8__b0_diff_11 = 0.0
+ sky130_fd_pr__pfet_01v8__b1_diff_11 = 0.0
+ sky130_fd_pr__pfet_01v8__agidl_diff_11 = 0.0
+ sky130_fd_pr__pfet_01v8__ua_diff_11 = -3.8915e-11
+ sky130_fd_pr__pfet_01v8__bgidl_diff_11 = 0.0
+ sky130_fd_pr__pfet_01v8__nfactor_diff_11 = 0.20363
+ sky130_fd_pr__pfet_01v8__ub_diff_11 = 4.9719e-19
+ sky130_fd_pr__pfet_01v8__pdits_diff_11 = 0.0
+ sky130_fd_pr__pfet_01v8__tvoff_diff_11 = 0.0
+ sky130_fd_pr__pfet_01v8__ags_diff_11 = 0.064145
+ sky130_fd_pr__pfet_01v8__k2_diff_11 = -0.014591
*
* sky130_fd_pr__pfet_01v8, Bin 012, W = 3.0, L = 2.0
* ---------------------------------
+ sky130_fd_pr__pfet_01v8__pdits_diff_12 = 0.0
+ sky130_fd_pr__pfet_01v8__tvoff_diff_12 = 0.0
+ sky130_fd_pr__pfet_01v8__ags_diff_12 = 0.05431
+ sky130_fd_pr__pfet_01v8__k2_diff_12 = -0.0081409
+ sky130_fd_pr__pfet_01v8__voff_diff_12 = -0.1031
+ sky130_fd_pr__pfet_01v8__a0_diff_12 = -0.060972
+ sky130_fd_pr__pfet_01v8__pditsd_diff_12 = 0.0
+ sky130_fd_pr__pfet_01v8__eta0_diff_12 = 0.0
+ sky130_fd_pr__pfet_01v8__vsat_diff_12 = 0.0
+ sky130_fd_pr__pfet_01v8__u0_diff_12 = 0.0024227
+ sky130_fd_pr__pfet_01v8__vth0_diff_12 = 0.0037563
+ sky130_fd_pr__pfet_01v8__cgidl_diff_12 = 0.0
+ sky130_fd_pr__pfet_01v8__keta_diff_12 = 0.0
+ sky130_fd_pr__pfet_01v8__rdsw_diff_12 = 0.0
+ sky130_fd_pr__pfet_01v8__kt1_diff_12 = 0.0
+ sky130_fd_pr__pfet_01v8__pclm_diff_12 = 0.0
+ sky130_fd_pr__pfet_01v8__b0_diff_12 = 0.0
+ sky130_fd_pr__pfet_01v8__b1_diff_12 = 0.0
+ sky130_fd_pr__pfet_01v8__agidl_diff_12 = 0.0
+ sky130_fd_pr__pfet_01v8__ua_diff_12 = -4.5581e-12
+ sky130_fd_pr__pfet_01v8__bgidl_diff_12 = 0.0
+ sky130_fd_pr__pfet_01v8__nfactor_diff_12 = 0.18632
+ sky130_fd_pr__pfet_01v8__ub_diff_12 = 5.4069e-19
*
* sky130_fd_pr__pfet_01v8, Bin 013, W = 3.0, L = 4.0
* ---------------------------------
+ sky130_fd_pr__pfet_01v8__bgidl_diff_13 = 0.0
+ sky130_fd_pr__pfet_01v8__nfactor_diff_13 = 0.18043
+ sky130_fd_pr__pfet_01v8__ub_diff_13 = 5.6615e-19
+ sky130_fd_pr__pfet_01v8__pdits_diff_13 = 0.0
+ sky130_fd_pr__pfet_01v8__tvoff_diff_13 = 0.0
+ sky130_fd_pr__pfet_01v8__ags_diff_13 = 0.020604
+ sky130_fd_pr__pfet_01v8__k2_diff_13 = -0.0062466
+ sky130_fd_pr__pfet_01v8__voff_diff_13 = -0.091816
+ sky130_fd_pr__pfet_01v8__a0_diff_13 = -0.023106
+ sky130_fd_pr__pfet_01v8__eta0_diff_13 = 0.0
+ sky130_fd_pr__pfet_01v8__pditsd_diff_13 = 0.0
+ sky130_fd_pr__pfet_01v8__u0_diff_13 = 0.002569
+ sky130_fd_pr__pfet_01v8__vsat_diff_13 = 0.0
+ sky130_fd_pr__pfet_01v8__vth0_diff_13 = 0.01316
+ sky130_fd_pr__pfet_01v8__cgidl_diff_13 = 0.0
+ sky130_fd_pr__pfet_01v8__keta_diff_13 = 0.0
+ sky130_fd_pr__pfet_01v8__rdsw_diff_13 = 0.0
+ sky130_fd_pr__pfet_01v8__kt1_diff_13 = 0.0
+ sky130_fd_pr__pfet_01v8__pclm_diff_13 = 0.0
+ sky130_fd_pr__pfet_01v8__b0_diff_13 = 0.0
+ sky130_fd_pr__pfet_01v8__b1_diff_13 = 0.0
+ sky130_fd_pr__pfet_01v8__agidl_diff_13 = 0.0
+ sky130_fd_pr__pfet_01v8__ua_diff_13 = -3.3779e-12
*
* sky130_fd_pr__pfet_01v8, Bin 014, W = 3.0, L = 8.0
* ---------------------------------
+ sky130_fd_pr__pfet_01v8__agidl_diff_14 = 0.0
+ sky130_fd_pr__pfet_01v8__b1_diff_14 = 0.0
+ sky130_fd_pr__pfet_01v8__ua_diff_14 = -3.0908e-12
+ sky130_fd_pr__pfet_01v8__bgidl_diff_14 = 0.0
+ sky130_fd_pr__pfet_01v8__nfactor_diff_14 = 0.20573
+ sky130_fd_pr__pfet_01v8__ub_diff_14 = 6.5948e-19
+ sky130_fd_pr__pfet_01v8__pdits_diff_14 = 0.0
+ sky130_fd_pr__pfet_01v8__tvoff_diff_14 = 0.0
+ sky130_fd_pr__pfet_01v8__ags_diff_14 = 0.0089123
+ sky130_fd_pr__pfet_01v8__k2_diff_14 = -0.0063904
+ sky130_fd_pr__pfet_01v8__voff_diff_14 = -0.083073
+ sky130_fd_pr__pfet_01v8__eta0_diff_14 = 0.0
+ sky130_fd_pr__pfet_01v8__a0_diff_14 = -0.010822
+ sky130_fd_pr__pfet_01v8__pditsd_diff_14 = 0.0
+ sky130_fd_pr__pfet_01v8__u0_diff_14 = 0.0030595
+ sky130_fd_pr__pfet_01v8__vsat_diff_14 = 0.0
+ sky130_fd_pr__pfet_01v8__vth0_diff_14 = 0.015683
+ sky130_fd_pr__pfet_01v8__cgidl_diff_14 = 0.0
+ sky130_fd_pr__pfet_01v8__keta_diff_14 = 0.0
+ sky130_fd_pr__pfet_01v8__rdsw_diff_14 = 0.0
+ sky130_fd_pr__pfet_01v8__kt1_diff_14 = 0.0
+ sky130_fd_pr__pfet_01v8__pclm_diff_14 = 0.0
+ sky130_fd_pr__pfet_01v8__b0_diff_14 = 0.0
*
* sky130_fd_pr__pfet_01v8, Bin 015, W = 3.0, L = 0.15
* ----------------------------------
+ sky130_fd_pr__pfet_01v8__b0_diff_15 = 0.0
+ sky130_fd_pr__pfet_01v8__agidl_diff_15 = 0.0
+ sky130_fd_pr__pfet_01v8__b1_diff_15 = 0.0
+ sky130_fd_pr__pfet_01v8__ua_diff_15 = 2.9356e-10
+ sky130_fd_pr__pfet_01v8__bgidl_diff_15 = 0.0
+ sky130_fd_pr__pfet_01v8__nfactor_diff_15 = 2.5923
+ sky130_fd_pr__pfet_01v8__ub_diff_15 = -5.5818e-20
+ sky130_fd_pr__pfet_01v8__tvoff_diff_15 = 0.0
+ sky130_fd_pr__pfet_01v8__ags_diff_15 = 0.0
+ sky130_fd_pr__pfet_01v8__k2_diff_15 = 0.00079783
+ sky130_fd_pr__pfet_01v8__pdits_diff_15 = 0.0
+ sky130_fd_pr__pfet_01v8__voff_diff_15 = -0.17313
+ sky130_fd_pr__pfet_01v8__eta0_diff_15 = 0.0
+ sky130_fd_pr__pfet_01v8__a0_diff_15 = 0.0
+ sky130_fd_pr__pfet_01v8__pditsd_diff_15 = 0.0
+ sky130_fd_pr__pfet_01v8__u0_diff_15 = 0.0011095
+ sky130_fd_pr__pfet_01v8__vsat_diff_15 = -20000.0
+ sky130_fd_pr__pfet_01v8__vth0_diff_15 = -0.16495
+ sky130_fd_pr__pfet_01v8__cgidl_diff_15 = 0.0
+ sky130_fd_pr__pfet_01v8__keta_diff_15 = 0.0
+ sky130_fd_pr__pfet_01v8__rdsw_diff_15 = 0.0
+ sky130_fd_pr__pfet_01v8__kt1_diff_15 = 0.0
+ sky130_fd_pr__pfet_01v8__pclm_diff_15 = 0.0
*
* sky130_fd_pr__pfet_01v8, Bin 016, W = 3.0, L = 0.18
* ----------------------------------
+ sky130_fd_pr__pfet_01v8__pclm_diff_16 = 0.0
+ sky130_fd_pr__pfet_01v8__b0_diff_16 = 0.0
+ sky130_fd_pr__pfet_01v8__agidl_diff_16 = 0.0
+ sky130_fd_pr__pfet_01v8__b1_diff_16 = 0.0
+ sky130_fd_pr__pfet_01v8__ua_diff_16 = 2.0851e-11
+ sky130_fd_pr__pfet_01v8__bgidl_diff_16 = 0.0
+ sky130_fd_pr__pfet_01v8__nfactor_diff_16 = 1.5107
+ sky130_fd_pr__pfet_01v8__tvoff_diff_16 = 0.0
+ sky130_fd_pr__pfet_01v8__ags_diff_16 = 0.0
+ sky130_fd_pr__pfet_01v8__ub_diff_16 = 1.946e-19
+ sky130_fd_pr__pfet_01v8__k2_diff_16 = 0.0030068
+ sky130_fd_pr__pfet_01v8__pdits_diff_16 = 0.0
+ sky130_fd_pr__pfet_01v8__voff_diff_16 = -0.27197
+ sky130_fd_pr__pfet_01v8__eta0_diff_16 = 0.0
+ sky130_fd_pr__pfet_01v8__a0_diff_16 = 0.0
+ sky130_fd_pr__pfet_01v8__pditsd_diff_16 = 0.0
+ sky130_fd_pr__pfet_01v8__u0_diff_16 = 0.00042752
+ sky130_fd_pr__pfet_01v8__vsat_diff_16 = -16788.0
+ sky130_fd_pr__pfet_01v8__vth0_diff_16 = -0.076492
+ sky130_fd_pr__pfet_01v8__cgidl_diff_16 = 0.0
+ sky130_fd_pr__pfet_01v8__keta_diff_16 = 0.0
+ sky130_fd_pr__pfet_01v8__rdsw_diff_16 = 0.0
+ sky130_fd_pr__pfet_01v8__kt1_diff_16 = 0.0
*
* sky130_fd_pr__pfet_01v8, Bin 017, W = 3.0, L = 0.25
* ----------------------------------
+ sky130_fd_pr__pfet_01v8__kt1_diff_17 = 0.0
+ sky130_fd_pr__pfet_01v8__pclm_diff_17 = 0.0
+ sky130_fd_pr__pfet_01v8__b0_diff_17 = 0.0
+ sky130_fd_pr__pfet_01v8__agidl_diff_17 = 0.0
+ sky130_fd_pr__pfet_01v8__b1_diff_17 = 0.0
+ sky130_fd_pr__pfet_01v8__bgidl_diff_17 = 0.0
+ sky130_fd_pr__pfet_01v8__nfactor_diff_17 = 0.83987
+ sky130_fd_pr__pfet_01v8__ua_diff_17 = -1.804e-11
+ sky130_fd_pr__pfet_01v8__tvoff_diff_17 = 0.0
+ sky130_fd_pr__pfet_01v8__ags_diff_17 = 0.0
+ sky130_fd_pr__pfet_01v8__ub_diff_17 = 2.52e-19
+ sky130_fd_pr__pfet_01v8__k2_diff_17 = 0.001971
+ sky130_fd_pr__pfet_01v8__pdits_diff_17 = 0.0
+ sky130_fd_pr__pfet_01v8__voff_diff_17 = -0.21242
+ sky130_fd_pr__pfet_01v8__eta0_diff_17 = 0.0
+ sky130_fd_pr__pfet_01v8__a0_diff_17 = 0.0
+ sky130_fd_pr__pfet_01v8__pditsd_diff_17 = 0.0
+ sky130_fd_pr__pfet_01v8__u0_diff_17 = 0.00027526
+ sky130_fd_pr__pfet_01v8__vsat_diff_17 = 30780.0
+ sky130_fd_pr__pfet_01v8__vth0_diff_17 = -0.031717
+ sky130_fd_pr__pfet_01v8__cgidl_diff_17 = 0.0
+ sky130_fd_pr__pfet_01v8__keta_diff_17 = 0.0
+ sky130_fd_pr__pfet_01v8__rdsw_diff_17 = 0.0
*
* sky130_fd_pr__pfet_01v8, Bin 018, W = 3.0, L = 0.5
* ---------------------------------
+ sky130_fd_pr__pfet_01v8__rdsw_diff_18 = 0.0
+ sky130_fd_pr__pfet_01v8__kt1_diff_18 = 0.0
+ sky130_fd_pr__pfet_01v8__pclm_diff_18 = 0.0
+ sky130_fd_pr__pfet_01v8__b0_diff_18 = 0.0
+ sky130_fd_pr__pfet_01v8__agidl_diff_18 = 0.0
+ sky130_fd_pr__pfet_01v8__b1_diff_18 = 0.0
+ sky130_fd_pr__pfet_01v8__bgidl_diff_18 = 0.0
+ sky130_fd_pr__pfet_01v8__nfactor_diff_18 = 0.51911
+ sky130_fd_pr__pfet_01v8__ua_diff_18 = 1.4339e-11
+ sky130_fd_pr__pfet_01v8__tvoff_diff_18 = 0.0
+ sky130_fd_pr__pfet_01v8__ags_diff_18 = 0.0
+ sky130_fd_pr__pfet_01v8__ub_diff_18 = 3.5515e-19
+ sky130_fd_pr__pfet_01v8__k2_diff_18 = -0.012538
+ sky130_fd_pr__pfet_01v8__pdits_diff_18 = 0.0
+ sky130_fd_pr__pfet_01v8__voff_diff_18 = -0.14187
+ sky130_fd_pr__pfet_01v8__eta0_diff_18 = 0.0
+ sky130_fd_pr__pfet_01v8__a0_diff_18 = 0.0
+ sky130_fd_pr__pfet_01v8__pditsd_diff_18 = 0.0
+ sky130_fd_pr__pfet_01v8__u0_diff_18 = 0.0013831
+ sky130_fd_pr__pfet_01v8__vsat_diff_18 = 15158.0
+ sky130_fd_pr__pfet_01v8__vth0_diff_18 = 0.01865
+ sky130_fd_pr__pfet_01v8__cgidl_diff_18 = 0.0
+ sky130_fd_pr__pfet_01v8__keta_diff_18 = 0.0
*
* sky130_fd_pr__pfet_01v8, Bin 019, W = 5.0, L = 1.0
* ---------------------------------
+ sky130_fd_pr__pfet_01v8__cgidl_diff_19 = 0.0
+ sky130_fd_pr__pfet_01v8__keta_diff_19 = 0.0
+ sky130_fd_pr__pfet_01v8__rdsw_diff_19 = 0.0
+ sky130_fd_pr__pfet_01v8__kt1_diff_19 = 0.0
+ sky130_fd_pr__pfet_01v8__pclm_diff_19 = 0.0
+ sky130_fd_pr__pfet_01v8__b0_diff_19 = 0.0
+ sky130_fd_pr__pfet_01v8__agidl_diff_19 = 0.0
+ sky130_fd_pr__pfet_01v8__b1_diff_19 = 0.0
+ sky130_fd_pr__pfet_01v8__bgidl_diff_19 = 0.0
+ sky130_fd_pr__pfet_01v8__nfactor_diff_19 = -0.041819
+ sky130_fd_pr__pfet_01v8__ua_diff_19 = -9.2578e-12
+ sky130_fd_pr__pfet_01v8__tvoff_diff_19 = 0.0
+ sky130_fd_pr__pfet_01v8__ags_diff_19 = 0.084095
+ sky130_fd_pr__pfet_01v8__ub_diff_19 = 3.6396e-19
+ sky130_fd_pr__pfet_01v8__k2_diff_19 = -0.009739
+ sky130_fd_pr__pfet_01v8__pdits_diff_19 = 0.0
+ sky130_fd_pr__pfet_01v8__voff_diff_19 = -0.091505
+ sky130_fd_pr__pfet_01v8__eta0_diff_19 = 0.0
+ sky130_fd_pr__pfet_01v8__a0_diff_19 = -0.084937
+ sky130_fd_pr__pfet_01v8__pditsd_diff_19 = 0.0
+ sky130_fd_pr__pfet_01v8__u0_diff_19 = 0.001464
+ sky130_fd_pr__pfet_01v8__vsat_diff_19 = 0.0
+ sky130_fd_pr__pfet_01v8__vth0_diff_19 = 0.021383
*
* sky130_fd_pr__pfet_01v8, Bin 020, W = 5.0, L = 2.0
* ---------------------------------
+ sky130_fd_pr__pfet_01v8__u0_diff_20 = 0.0016533
+ sky130_fd_pr__pfet_01v8__vth0_diff_20 = 0.016618
+ sky130_fd_pr__pfet_01v8__cgidl_diff_20 = 0.0
+ sky130_fd_pr__pfet_01v8__keta_diff_20 = 0.0
+ sky130_fd_pr__pfet_01v8__rdsw_diff_20 = 0.0
+ sky130_fd_pr__pfet_01v8__kt1_diff_20 = 0.0
+ sky130_fd_pr__pfet_01v8__pclm_diff_20 = 0.0
+ sky130_fd_pr__pfet_01v8__b0_diff_20 = 0.0
+ sky130_fd_pr__pfet_01v8__b1_diff_20 = 0.0
+ sky130_fd_pr__pfet_01v8__agidl_diff_20 = 0.0
+ sky130_fd_pr__pfet_01v8__ua_diff_20 = -2.3869e-12
+ sky130_fd_pr__pfet_01v8__bgidl_diff_20 = 0.0
+ sky130_fd_pr__pfet_01v8__nfactor_diff_20 = 0.19236
+ sky130_fd_pr__pfet_01v8__ub_diff_20 = 3.5988e-19
+ sky130_fd_pr__pfet_01v8__pdits_diff_20 = 0.0
+ sky130_fd_pr__pfet_01v8__tvoff_diff_20 = 0.0
+ sky130_fd_pr__pfet_01v8__ags_diff_20 = 0.010814
+ sky130_fd_pr__pfet_01v8__k2_diff_20 = -0.0091133
+ sky130_fd_pr__pfet_01v8__voff_diff_20 = -0.085869
+ sky130_fd_pr__pfet_01v8__a0_diff_20 = -0.011877
+ sky130_fd_pr__pfet_01v8__pditsd_diff_20 = 0.0
+ sky130_fd_pr__pfet_01v8__eta0_diff_20 = 0.0
+ sky130_fd_pr__pfet_01v8__vsat_diff_20 = 0.0
*
* sky130_fd_pr__pfet_01v8, Bin 021, W = 5.0, L = 4.0
* ---------------------------------
+ sky130_fd_pr__pfet_01v8__pditsd_diff_21 = 0.0
+ sky130_fd_pr__pfet_01v8__eta0_diff_21 = 0.0
+ sky130_fd_pr__pfet_01v8__vsat_diff_21 = 0.0
+ sky130_fd_pr__pfet_01v8__u0_diff_21 = 0.0022548
+ sky130_fd_pr__pfet_01v8__vth0_diff_21 = 0.019913
+ sky130_fd_pr__pfet_01v8__cgidl_diff_21 = 0.0
+ sky130_fd_pr__pfet_01v8__keta_diff_21 = 0.0
+ sky130_fd_pr__pfet_01v8__rdsw_diff_21 = 0.0
+ sky130_fd_pr__pfet_01v8__kt1_diff_21 = 0.0
+ sky130_fd_pr__pfet_01v8__pclm_diff_21 = 0.0
+ sky130_fd_pr__pfet_01v8__b0_diff_21 = 0.0
+ sky130_fd_pr__pfet_01v8__b1_diff_21 = 0.0
+ sky130_fd_pr__pfet_01v8__agidl_diff_21 = 0.0
+ sky130_fd_pr__pfet_01v8__ua_diff_21 = -4.1623e-12
+ sky130_fd_pr__pfet_01v8__bgidl_diff_21 = 0.0
+ sky130_fd_pr__pfet_01v8__nfactor_diff_21 = 0.14933
+ sky130_fd_pr__pfet_01v8__ub_diff_21 = 4.7009e-19
+ sky130_fd_pr__pfet_01v8__pdits_diff_21 = 0.0
+ sky130_fd_pr__pfet_01v8__tvoff_diff_21 = 0.0
+ sky130_fd_pr__pfet_01v8__ags_diff_21 = 0.0073418
+ sky130_fd_pr__pfet_01v8__k2_diff_21 = -0.0096588
+ sky130_fd_pr__pfet_01v8__voff_diff_21 = -0.081178
+ sky130_fd_pr__pfet_01v8__a0_diff_21 = -0.0082007
*
* sky130_fd_pr__pfet_01v8, Bin 022, W = 5.0, L = 8.0
* ---------------------------------
+ sky130_fd_pr__pfet_01v8__voff_diff_22 = -0.078696
+ sky130_fd_pr__pfet_01v8__a0_diff_22 = -0.011308
+ sky130_fd_pr__pfet_01v8__pditsd_diff_22 = 0.0
+ sky130_fd_pr__pfet_01v8__eta0_diff_22 = 0.0
+ sky130_fd_pr__pfet_01v8__vsat_diff_22 = 0.0
+ sky130_fd_pr__pfet_01v8__u0_diff_22 = 0.00247
+ sky130_fd_pr__pfet_01v8__vth0_diff_22 = 0.013766
+ sky130_fd_pr__pfet_01v8__cgidl_diff_22 = 0.0
+ sky130_fd_pr__pfet_01v8__keta_diff_22 = 0.0
+ sky130_fd_pr__pfet_01v8__rdsw_diff_22 = 0.0
+ sky130_fd_pr__pfet_01v8__kt1_diff_22 = 0.0
+ sky130_fd_pr__pfet_01v8__pclm_diff_22 = 0.0
+ sky130_fd_pr__pfet_01v8__b0_diff_22 = 0.0
+ sky130_fd_pr__pfet_01v8__b1_diff_22 = 0.0
+ sky130_fd_pr__pfet_01v8__agidl_diff_22 = 0.0
+ sky130_fd_pr__pfet_01v8__ua_diff_22 = -2.2073e-12
+ sky130_fd_pr__pfet_01v8__bgidl_diff_22 = 0.0
+ sky130_fd_pr__pfet_01v8__nfactor_diff_22 = 0.21399
+ sky130_fd_pr__pfet_01v8__ub_diff_22 = 5.0422e-19
+ sky130_fd_pr__pfet_01v8__pdits_diff_22 = 0.0
+ sky130_fd_pr__pfet_01v8__tvoff_diff_22 = 0.0
+ sky130_fd_pr__pfet_01v8__ags_diff_22 = 0.010315
+ sky130_fd_pr__pfet_01v8__k2_diff_22 = -0.009782
*
* sky130_fd_pr__pfet_01v8, Bin 023, W = 5.0, L = 0.15
* ----------------------------------
+ sky130_fd_pr__pfet_01v8__pdits_diff_23 = 0.0
+ sky130_fd_pr__pfet_01v8__tvoff_diff_23 = 0.0
+ sky130_fd_pr__pfet_01v8__ags_diff_23 = 0.0
+ sky130_fd_pr__pfet_01v8__k2_diff_23 = 0.040345
+ sky130_fd_pr__pfet_01v8__voff_diff_23 = -0.16849
+ sky130_fd_pr__pfet_01v8__a0_diff_23 = 0.0
+ sky130_fd_pr__pfet_01v8__pditsd_diff_23 = 0.0
+ sky130_fd_pr__pfet_01v8__eta0_diff_23 = 0.0
+ sky130_fd_pr__pfet_01v8__vsat_diff_23 = -20000.0
+ sky130_fd_pr__pfet_01v8__u0_diff_23 = -0.001202
+ sky130_fd_pr__pfet_01v8__vth0_diff_23 = -0.095482
+ sky130_fd_pr__pfet_01v8__cgidl_diff_23 = 0.0
+ sky130_fd_pr__pfet_01v8__keta_diff_23 = 0.0
+ sky130_fd_pr__pfet_01v8__rdsw_diff_23 = 0.0
+ sky130_fd_pr__pfet_01v8__kt1_diff_23 = 0.0
+ sky130_fd_pr__pfet_01v8__pclm_diff_23 = 0.0
+ sky130_fd_pr__pfet_01v8__b0_diff_23 = 0.0
+ sky130_fd_pr__pfet_01v8__b1_diff_23 = 0.0
+ sky130_fd_pr__pfet_01v8__agidl_diff_23 = 0.0
+ sky130_fd_pr__pfet_01v8__ua_diff_23 = -4.5385e-10
+ sky130_fd_pr__pfet_01v8__bgidl_diff_23 = 0.0
+ sky130_fd_pr__pfet_01v8__nfactor_diff_23 = 1.3313
+ sky130_fd_pr__pfet_01v8__ub_diff_23 = 4.7501e-19
*
* sky130_fd_pr__pfet_01v8, Bin 024, W = 5.0, L = 0.18
* ----------------------------------
+ sky130_fd_pr__pfet_01v8__bgidl_diff_24 = 0.0
+ sky130_fd_pr__pfet_01v8__nfactor_diff_24 = 1.5511
+ sky130_fd_pr__pfet_01v8__ub_diff_24 = 1.4305e-19
+ sky130_fd_pr__pfet_01v8__pdits_diff_24 = 0.0
+ sky130_fd_pr__pfet_01v8__tvoff_diff_24 = 0.0
+ sky130_fd_pr__pfet_01v8__ags_diff_24 = 0.0
+ sky130_fd_pr__pfet_01v8__k2_diff_24 = 0.0052883
+ sky130_fd_pr__pfet_01v8__voff_diff_24 = -0.25463
+ sky130_fd_pr__pfet_01v8__a0_diff_24 = 0.0
+ sky130_fd_pr__pfet_01v8__eta0_diff_24 = 0.0
+ sky130_fd_pr__pfet_01v8__pditsd_diff_24 = 0.0
+ sky130_fd_pr__pfet_01v8__u0_diff_24 = 9.8714e-5
+ sky130_fd_pr__pfet_01v8__vsat_diff_24 = -3689.3
+ sky130_fd_pr__pfet_01v8__vth0_diff_24 = -0.090211
+ sky130_fd_pr__pfet_01v8__cgidl_diff_24 = 0.0
+ sky130_fd_pr__pfet_01v8__keta_diff_24 = 0.0
+ sky130_fd_pr__pfet_01v8__rdsw_diff_24 = 0.0
+ sky130_fd_pr__pfet_01v8__kt1_diff_24 = 0.0
+ sky130_fd_pr__pfet_01v8__pclm_diff_24 = 0.0
+ sky130_fd_pr__pfet_01v8__b0_diff_24 = 0.0
+ sky130_fd_pr__pfet_01v8__b1_diff_24 = 0.0
+ sky130_fd_pr__pfet_01v8__agidl_diff_24 = 0.0
+ sky130_fd_pr__pfet_01v8__ua_diff_24 = -5.787e-12
*
* sky130_fd_pr__pfet_01v8, Bin 025, W = 5.0, L = 0.25
* ----------------------------------
+ sky130_fd_pr__pfet_01v8__agidl_diff_25 = 0.0
+ sky130_fd_pr__pfet_01v8__b1_diff_25 = 0.0
+ sky130_fd_pr__pfet_01v8__ua_diff_25 = 1.5952e-12
+ sky130_fd_pr__pfet_01v8__bgidl_diff_25 = 0.0
+ sky130_fd_pr__pfet_01v8__nfactor_diff_25 = 0.56131
+ sky130_fd_pr__pfet_01v8__ub_diff_25 = 2.0125e-19
+ sky130_fd_pr__pfet_01v8__pdits_diff_25 = 0.0
+ sky130_fd_pr__pfet_01v8__tvoff_diff_25 = 0.0
+ sky130_fd_pr__pfet_01v8__ags_diff_25 = 0.0
+ sky130_fd_pr__pfet_01v8__k2_diff_25 = -0.00017766
+ sky130_fd_pr__pfet_01v8__voff_diff_25 = -0.20387
+ sky130_fd_pr__pfet_01v8__eta0_diff_25 = 0.0
+ sky130_fd_pr__pfet_01v8__a0_diff_25 = 0.0
+ sky130_fd_pr__pfet_01v8__pditsd_diff_25 = 0.0
+ sky130_fd_pr__pfet_01v8__u0_diff_25 = 0.00043733
+ sky130_fd_pr__pfet_01v8__vsat_diff_25 = 4289.2
+ sky130_fd_pr__pfet_01v8__vth0_diff_25 = -0.0463
+ sky130_fd_pr__pfet_01v8__cgidl_diff_25 = 0.0
+ sky130_fd_pr__pfet_01v8__keta_diff_25 = 0.0
+ sky130_fd_pr__pfet_01v8__rdsw_diff_25 = 0.0
+ sky130_fd_pr__pfet_01v8__kt1_diff_25 = 0.0
+ sky130_fd_pr__pfet_01v8__pclm_diff_25 = 0.0
+ sky130_fd_pr__pfet_01v8__b0_diff_25 = 0.0
*
* sky130_fd_pr__pfet_01v8, Bin 026, W = 5.0, L = 0.5
* ---------------------------------
+ sky130_fd_pr__pfet_01v8__b0_diff_26 = 0.0
+ sky130_fd_pr__pfet_01v8__agidl_diff_26 = 0.0
+ sky130_fd_pr__pfet_01v8__b1_diff_26 = 0.0
+ sky130_fd_pr__pfet_01v8__ua_diff_26 = 2.4056e-11
+ sky130_fd_pr__pfet_01v8__bgidl_diff_26 = 0.0
+ sky130_fd_pr__pfet_01v8__nfactor_diff_26 = 0.3907
+ sky130_fd_pr__pfet_01v8__ub_diff_26 = 3.3049e-19
+ sky130_fd_pr__pfet_01v8__tvoff_diff_26 = 0.0
+ sky130_fd_pr__pfet_01v8__ags_diff_26 = 0.0
+ sky130_fd_pr__pfet_01v8__k2_diff_26 = -0.011709
+ sky130_fd_pr__pfet_01v8__pdits_diff_26 = 0.0
+ sky130_fd_pr__pfet_01v8__voff_diff_26 = -0.098432
+ sky130_fd_pr__pfet_01v8__eta0_diff_26 = 0.0
+ sky130_fd_pr__pfet_01v8__a0_diff_26 = 0.0
+ sky130_fd_pr__pfet_01v8__pditsd_diff_26 = 0.0
+ sky130_fd_pr__pfet_01v8__u0_diff_26 = 0.0015274
+ sky130_fd_pr__pfet_01v8__vsat_diff_26 = -7322.9
+ sky130_fd_pr__pfet_01v8__vth0_diff_26 = 0.01124
+ sky130_fd_pr__pfet_01v8__cgidl_diff_26 = 0.0
+ sky130_fd_pr__pfet_01v8__keta_diff_26 = 0.0
+ sky130_fd_pr__pfet_01v8__rdsw_diff_26 = 0.0
+ sky130_fd_pr__pfet_01v8__kt1_diff_26 = 0.0
+ sky130_fd_pr__pfet_01v8__pclm_diff_26 = 0.0
*
* sky130_fd_pr__pfet_01v8, Bin 027, W = 7.0, L = 1.0
* ---------------------------------
+ sky130_fd_pr__pfet_01v8__pclm_diff_27 = 0.0
+ sky130_fd_pr__pfet_01v8__b0_diff_27 = 0.0
+ sky130_fd_pr__pfet_01v8__agidl_diff_27 = 0.0
+ sky130_fd_pr__pfet_01v8__b1_diff_27 = 0.0
+ sky130_fd_pr__pfet_01v8__ua_diff_27 = 6.4042e-12
+ sky130_fd_pr__pfet_01v8__bgidl_diff_27 = 0.0
+ sky130_fd_pr__pfet_01v8__nfactor_diff_27 = 0.039245
+ sky130_fd_pr__pfet_01v8__tvoff_diff_27 = 0.0
+ sky130_fd_pr__pfet_01v8__ags_diff_27 = 0.083559
+ sky130_fd_pr__pfet_01v8__ub_diff_27 = 3.8976e-19
+ sky130_fd_pr__pfet_01v8__k2_diff_27 = -0.0083062
+ sky130_fd_pr__pfet_01v8__pdits_diff_27 = 0.0
+ sky130_fd_pr__pfet_01v8__voff_diff_27 = -0.072852
+ sky130_fd_pr__pfet_01v8__eta0_diff_27 = 0.0
+ sky130_fd_pr__pfet_01v8__a0_diff_27 = -0.11904
+ sky130_fd_pr__pfet_01v8__pditsd_diff_27 = 0.0
+ sky130_fd_pr__pfet_01v8__u0_diff_27 = 0.0017166
+ sky130_fd_pr__pfet_01v8__vsat_diff_27 = 0.0
+ sky130_fd_pr__pfet_01v8__vth0_diff_27 = 0.010829
+ sky130_fd_pr__pfet_01v8__cgidl_diff_27 = 0.0
+ sky130_fd_pr__pfet_01v8__keta_diff_27 = 0.0
+ sky130_fd_pr__pfet_01v8__rdsw_diff_27 = 0.0
+ sky130_fd_pr__pfet_01v8__kt1_diff_27 = 0.0
*
* sky130_fd_pr__pfet_01v8, Bin 028, W = 7.0, L = 2.0
* ---------------------------------
+ sky130_fd_pr__pfet_01v8__kt1_diff_28 = 0.0
+ sky130_fd_pr__pfet_01v8__pclm_diff_28 = 0.0
+ sky130_fd_pr__pfet_01v8__b0_diff_28 = 0.0
+ sky130_fd_pr__pfet_01v8__agidl_diff_28 = 0.0
+ sky130_fd_pr__pfet_01v8__b1_diff_28 = 0.0
+ sky130_fd_pr__pfet_01v8__bgidl_diff_28 = 0.0
+ sky130_fd_pr__pfet_01v8__nfactor_diff_28 = 0.10842
+ sky130_fd_pr__pfet_01v8__ua_diff_28 = -3.7462e-12
+ sky130_fd_pr__pfet_01v8__tvoff_diff_28 = 0.0
+ sky130_fd_pr__pfet_01v8__ags_diff_28 = 0.055844
+ sky130_fd_pr__pfet_01v8__ub_diff_28 = 3.9115e-19
+ sky130_fd_pr__pfet_01v8__k2_diff_28 = -0.010797
+ sky130_fd_pr__pfet_01v8__pdits_diff_28 = 0.0
+ sky130_fd_pr__pfet_01v8__voff_diff_28 = -0.078111
+ sky130_fd_pr__pfet_01v8__eta0_diff_28 = 0.0
+ sky130_fd_pr__pfet_01v8__a0_diff_28 = -0.061503
+ sky130_fd_pr__pfet_01v8__pditsd_diff_28 = 0.0
+ sky130_fd_pr__pfet_01v8__u0_diff_28 = 0.0018235
+ sky130_fd_pr__pfet_01v8__vsat_diff_28 = 0.0
+ sky130_fd_pr__pfet_01v8__vth0_diff_28 = 0.018136
+ sky130_fd_pr__pfet_01v8__cgidl_diff_28 = 0.0
+ sky130_fd_pr__pfet_01v8__keta_diff_28 = 0.0
+ sky130_fd_pr__pfet_01v8__rdsw_diff_28 = 0.0
*
* sky130_fd_pr__pfet_01v8, Bin 029, W = 7.0, L = 4.0
* ---------------------------------
+ sky130_fd_pr__pfet_01v8__rdsw_diff_29 = 0.0
+ sky130_fd_pr__pfet_01v8__kt1_diff_29 = 0.0
+ sky130_fd_pr__pfet_01v8__pclm_diff_29 = 0.0
+ sky130_fd_pr__pfet_01v8__b0_diff_29 = 0.0
+ sky130_fd_pr__pfet_01v8__agidl_diff_29 = 0.0
+ sky130_fd_pr__pfet_01v8__b1_diff_29 = 0.0
+ sky130_fd_pr__pfet_01v8__bgidl_diff_29 = 0.0
+ sky130_fd_pr__pfet_01v8__nfactor_diff_29 = 0.18611
+ sky130_fd_pr__pfet_01v8__ua_diff_29 = -1.9042e-12
+ sky130_fd_pr__pfet_01v8__tvoff_diff_29 = 0.0
+ sky130_fd_pr__pfet_01v8__ags_diff_29 = 0.014379
+ sky130_fd_pr__pfet_01v8__ub_diff_29 = 5.042e-19
+ sky130_fd_pr__pfet_01v8__k2_diff_29 = -0.010381
+ sky130_fd_pr__pfet_01v8__pdits_diff_29 = 0.0
+ sky130_fd_pr__pfet_01v8__voff_diff_29 = -0.0803
+ sky130_fd_pr__pfet_01v8__eta0_diff_29 = 0.0
+ sky130_fd_pr__pfet_01v8__a0_diff_29 = -0.017759
+ sky130_fd_pr__pfet_01v8__pditsd_diff_29 = 0.0
+ sky130_fd_pr__pfet_01v8__u0_diff_29 = 0.0025177
+ sky130_fd_pr__pfet_01v8__vsat_diff_29 = 0.0
+ sky130_fd_pr__pfet_01v8__vth0_diff_29 = 0.013702
+ sky130_fd_pr__pfet_01v8__cgidl_diff_29 = 0.0
+ sky130_fd_pr__pfet_01v8__keta_diff_29 = 0.0
*
* sky130_fd_pr__pfet_01v8, Bin 030, W = 7.0, L = 8.0
* ---------------------------------
+ sky130_fd_pr__pfet_01v8__cgidl_diff_30 = 0.0
+ sky130_fd_pr__pfet_01v8__keta_diff_30 = 0.0
+ sky130_fd_pr__pfet_01v8__rdsw_diff_30 = 0.0
+ sky130_fd_pr__pfet_01v8__kt1_diff_30 = 0.0
+ sky130_fd_pr__pfet_01v8__pclm_diff_30 = 0.0
+ sky130_fd_pr__pfet_01v8__b0_diff_30 = 0.0
+ sky130_fd_pr__pfet_01v8__b1_diff_30 = 0.0
+ sky130_fd_pr__pfet_01v8__agidl_diff_30 = 0.0
+ sky130_fd_pr__pfet_01v8__ua_diff_30 = -5.5272e-12
+ sky130_fd_pr__pfet_01v8__bgidl_diff_30 = 0.0
+ sky130_fd_pr__pfet_01v8__nfactor_diff_30 = 0.28527
+ sky130_fd_pr__pfet_01v8__ub_diff_30 = 5.2353e-19
+ sky130_fd_pr__pfet_01v8__pdits_diff_30 = 0.0
+ sky130_fd_pr__pfet_01v8__tvoff_diff_30 = 0.0
+ sky130_fd_pr__pfet_01v8__ags_diff_30 = 0.020428
+ sky130_fd_pr__pfet_01v8__k2_diff_30 = -0.010828
+ sky130_fd_pr__pfet_01v8__voff_diff_30 = -0.088406
+ sky130_fd_pr__pfet_01v8__a0_diff_30 = -0.021977
+ sky130_fd_pr__pfet_01v8__pditsd_diff_30 = 0.0
+ sky130_fd_pr__pfet_01v8__eta0_diff_30 = 0.0
+ sky130_fd_pr__pfet_01v8__vsat_diff_30 = 0.0
+ sky130_fd_pr__pfet_01v8__u0_diff_30 = 0.0026341
+ sky130_fd_pr__pfet_01v8__vth0_diff_30 = 0.011346
*
* sky130_fd_pr__pfet_01v8, Bin 031, W = 7.0, L = 0.15
* ----------------------------------
+ sky130_fd_pr__pfet_01v8__u0_diff_31 = 3.7129e-5
+ sky130_fd_pr__pfet_01v8__vth0_diff_31 = -0.15789
+ sky130_fd_pr__pfet_01v8__cgidl_diff_31 = 0.0
+ sky130_fd_pr__pfet_01v8__keta_diff_31 = 0.0
+ sky130_fd_pr__pfet_01v8__rdsw_diff_31 = 0.0
+ sky130_fd_pr__pfet_01v8__kt1_diff_31 = 0.0
+ sky130_fd_pr__pfet_01v8__pclm_diff_31 = 0.0
+ sky130_fd_pr__pfet_01v8__b0_diff_31 = 0.0
+ sky130_fd_pr__pfet_01v8__b1_diff_31 = 0.0
+ sky130_fd_pr__pfet_01v8__agidl_diff_31 = 0.0
+ sky130_fd_pr__pfet_01v8__ua_diff_31 = -2.4799e-11
+ sky130_fd_pr__pfet_01v8__bgidl_diff_31 = 0.0
+ sky130_fd_pr__pfet_01v8__nfactor_diff_31 = 1.7187
+ sky130_fd_pr__pfet_01v8__ub_diff_31 = 1.2123e-19
+ sky130_fd_pr__pfet_01v8__pdits_diff_31 = 0.0
+ sky130_fd_pr__pfet_01v8__tvoff_diff_31 = 0.0
+ sky130_fd_pr__pfet_01v8__ags_diff_31 = 0.0
+ sky130_fd_pr__pfet_01v8__k2_diff_31 = 0.0033879
+ sky130_fd_pr__pfet_01v8__voff_diff_31 = -0.19076
+ sky130_fd_pr__pfet_01v8__a0_diff_31 = 0.0
+ sky130_fd_pr__pfet_01v8__pditsd_diff_31 = 0.0
+ sky130_fd_pr__pfet_01v8__eta0_diff_31 = 0.0
+ sky130_fd_pr__pfet_01v8__vsat_diff_31 = -16802.0
*
* sky130_fd_pr__pfet_01v8, Bin 032, W = 7.0, L = 0.18
* ----------------------------------
+ sky130_fd_pr__pfet_01v8__pditsd_diff_32 = 0.0
+ sky130_fd_pr__pfet_01v8__eta0_diff_32 = 0.0
+ sky130_fd_pr__pfet_01v8__vsat_diff_32 = -8920.3
+ sky130_fd_pr__pfet_01v8__u0_diff_32 = 0.00019198
+ sky130_fd_pr__pfet_01v8__vth0_diff_32 = -0.091404
+ sky130_fd_pr__pfet_01v8__cgidl_diff_32 = 0.0
+ sky130_fd_pr__pfet_01v8__keta_diff_32 = 0.0
+ sky130_fd_pr__pfet_01v8__rdsw_diff_32 = 0.0
+ sky130_fd_pr__pfet_01v8__kt1_diff_32 = 0.0
+ sky130_fd_pr__pfet_01v8__pclm_diff_32 = 0.0
+ sky130_fd_pr__pfet_01v8__b0_diff_32 = 0.0
+ sky130_fd_pr__pfet_01v8__b1_diff_32 = 0.0
+ sky130_fd_pr__pfet_01v8__agidl_diff_32 = 0.0
+ sky130_fd_pr__pfet_01v8__ua_diff_32 = 1.8792e-11
+ sky130_fd_pr__pfet_01v8__bgidl_diff_32 = 0.0
+ sky130_fd_pr__pfet_01v8__nfactor_diff_32 = 0.97661
+ sky130_fd_pr__pfet_01v8__ub_diff_32 = 1.0728e-19
+ sky130_fd_pr__pfet_01v8__pdits_diff_32 = 0.0
+ sky130_fd_pr__pfet_01v8__tvoff_diff_32 = 0.0
+ sky130_fd_pr__pfet_01v8__ags_diff_32 = 0.0
+ sky130_fd_pr__pfet_01v8__k2_diff_32 = 0.0012343
+ sky130_fd_pr__pfet_01v8__voff_diff_32 = -0.16126
+ sky130_fd_pr__pfet_01v8__a0_diff_32 = 0.0
*
* sky130_fd_pr__pfet_01v8, Bin 033, W = 7.0, L = 0.25
* ----------------------------------
+ sky130_fd_pr__pfet_01v8__voff_diff_33 = -0.13694
+ sky130_fd_pr__pfet_01v8__a0_diff_33 = 0.0
+ sky130_fd_pr__pfet_01v8__pditsd_diff_33 = 0.0
+ sky130_fd_pr__pfet_01v8__eta0_diff_33 = 0.0
+ sky130_fd_pr__pfet_01v8__vsat_diff_33 = 8184.4
+ sky130_fd_pr__pfet_01v8__u0_diff_33 = 0.00037449
+ sky130_fd_pr__pfet_01v8__vth0_diff_33 = -0.043302
+ sky130_fd_pr__pfet_01v8__cgidl_diff_33 = 0.0
+ sky130_fd_pr__pfet_01v8__keta_diff_33 = 0.0
+ sky130_fd_pr__pfet_01v8__rdsw_diff_33 = 0.0
+ sky130_fd_pr__pfet_01v8__kt1_diff_33 = 0.0
+ sky130_fd_pr__pfet_01v8__pclm_diff_33 = 0.0
+ sky130_fd_pr__pfet_01v8__b0_diff_33 = 0.0
+ sky130_fd_pr__pfet_01v8__b1_diff_33 = 0.0
+ sky130_fd_pr__pfet_01v8__agidl_diff_33 = 0.0
+ sky130_fd_pr__pfet_01v8__ua_diff_33 = 3.1868e-12
+ sky130_fd_pr__pfet_01v8__bgidl_diff_33 = 0.0
+ sky130_fd_pr__pfet_01v8__nfactor_diff_33 = 0.32299
+ sky130_fd_pr__pfet_01v8__ub_diff_33 = 1.7315e-19
+ sky130_fd_pr__pfet_01v8__pdits_diff_33 = 0.0
+ sky130_fd_pr__pfet_01v8__tvoff_diff_33 = 0.0
+ sky130_fd_pr__pfet_01v8__ags_diff_33 = 0.0
+ sky130_fd_pr__pfet_01v8__k2_diff_33 = -0.0032062
*
* sky130_fd_pr__pfet_01v8, Bin 034, W = 7.0, L = 0.5
* ---------------------------------
+ sky130_fd_pr__pfet_01v8__pdits_diff_34 = 0.0
+ sky130_fd_pr__pfet_01v8__tvoff_diff_34 = 0.0
+ sky130_fd_pr__pfet_01v8__ags_diff_34 = 0.0
+ sky130_fd_pr__pfet_01v8__k2_diff_34 = -0.014635
+ sky130_fd_pr__pfet_01v8__voff_diff_34 = -0.10994
+ sky130_fd_pr__pfet_01v8__a0_diff_34 = 0.0
+ sky130_fd_pr__pfet_01v8__pditsd_diff_34 = 0.0
+ sky130_fd_pr__pfet_01v8__eta0_diff_34 = 0.0
+ sky130_fd_pr__pfet_01v8__vsat_diff_34 = 18609.0
+ sky130_fd_pr__pfet_01v8__u0_diff_34 = 0.0015571
+ sky130_fd_pr__pfet_01v8__vth0_diff_34 = -0.0010985
+ sky130_fd_pr__pfet_01v8__cgidl_diff_34 = 0.0
+ sky130_fd_pr__pfet_01v8__keta_diff_34 = 0.0
+ sky130_fd_pr__pfet_01v8__rdsw_diff_34 = 0.0
+ sky130_fd_pr__pfet_01v8__kt1_diff_34 = 0.0
+ sky130_fd_pr__pfet_01v8__pclm_diff_34 = 0.0
+ sky130_fd_pr__pfet_01v8__b0_diff_34 = 0.0
+ sky130_fd_pr__pfet_01v8__b1_diff_34 = 0.0
+ sky130_fd_pr__pfet_01v8__agidl_diff_34 = 0.0
+ sky130_fd_pr__pfet_01v8__ua_diff_34 = 3.2727e-12
+ sky130_fd_pr__pfet_01v8__bgidl_diff_34 = 0.0
+ sky130_fd_pr__pfet_01v8__nfactor_diff_34 = 0.24718
+ sky130_fd_pr__pfet_01v8__ub_diff_34 = 3.9575e-19
*
* sky130_fd_pr__pfet_01v8, Bin 035, W = 0.42, L = 1.0
* ----------------------------------
+ sky130_fd_pr__pfet_01v8__bgidl_diff_35 = 0.0
+ sky130_fd_pr__pfet_01v8__nfactor_diff_35 = 0.90855
+ sky130_fd_pr__pfet_01v8__ub_diff_35 = 6.0253e-19
+ sky130_fd_pr__pfet_01v8__pdits_diff_35 = 0.0
+ sky130_fd_pr__pfet_01v8__tvoff_diff_35 = 0.0
+ sky130_fd_pr__pfet_01v8__ags_diff_35 = 0.0
+ sky130_fd_pr__pfet_01v8__k2_diff_35 = -0.0086286
+ sky130_fd_pr__pfet_01v8__voff_diff_35 = -0.18543
+ sky130_fd_pr__pfet_01v8__a0_diff_35 = 0.0
+ sky130_fd_pr__pfet_01v8__eta0_diff_35 = 0.0
+ sky130_fd_pr__pfet_01v8__pditsd_diff_35 = 0.0
+ sky130_fd_pr__pfet_01v8__u0_diff_35 = 0.002693
+ sky130_fd_pr__pfet_01v8__vsat_diff_35 = 0.0
+ sky130_fd_pr__pfet_01v8__vth0_diff_35 = 0.013624
+ sky130_fd_pr__pfet_01v8__cgidl_diff_35 = 0.0
+ sky130_fd_pr__pfet_01v8__keta_diff_35 = 0.0
+ sky130_fd_pr__pfet_01v8__rdsw_diff_35 = 0.0
+ sky130_fd_pr__pfet_01v8__kt1_diff_35 = 0.0
+ sky130_fd_pr__pfet_01v8__pclm_diff_35 = 0.0
+ sky130_fd_pr__pfet_01v8__b0_diff_35 = 1.3259e-8
+ sky130_fd_pr__pfet_01v8__b1_diff_35 = 1.0302e-8
+ sky130_fd_pr__pfet_01v8__agidl_diff_35 = 0.0
+ sky130_fd_pr__pfet_01v8__ua_diff_35 = 1.3766e-12
*
* sky130_fd_pr__pfet_01v8, Bin 036, W = 0.42, L = 20.0
* -----------------------------------
+ sky130_fd_pr__pfet_01v8__agidl_diff_36 = 0.0
+ sky130_fd_pr__pfet_01v8__b1_diff_36 = 2.4775e-9
+ sky130_fd_pr__pfet_01v8__ua_diff_36 = -3.2012e-11
+ sky130_fd_pr__pfet_01v8__bgidl_diff_36 = 0.0
+ sky130_fd_pr__pfet_01v8__nfactor_diff_36 = 0.59531
+ sky130_fd_pr__pfet_01v8__ub_diff_36 = 2.0645e-20
+ sky130_fd_pr__pfet_01v8__pdits_diff_36 = 0.0
+ sky130_fd_pr__pfet_01v8__tvoff_diff_36 = 0.0
+ sky130_fd_pr__pfet_01v8__ags_diff_36 = 0.0
+ sky130_fd_pr__pfet_01v8__k2_diff_36 = -0.0021702
+ sky130_fd_pr__pfet_01v8__voff_diff_36 = -0.11002
+ sky130_fd_pr__pfet_01v8__eta0_diff_36 = 0.0
+ sky130_fd_pr__pfet_01v8__a0_diff_36 = 0.0
+ sky130_fd_pr__pfet_01v8__pditsd_diff_36 = 0.0
+ sky130_fd_pr__pfet_01v8__u0_diff_36 = -0.00028449
+ sky130_fd_pr__pfet_01v8__vsat_diff_36 = 20006.0
+ sky130_fd_pr__pfet_01v8__vth0_diff_36 = 0.036132
+ sky130_fd_pr__pfet_01v8__cgidl_diff_36 = 0.0
+ sky130_fd_pr__pfet_01v8__keta_diff_36 = 0.0
+ sky130_fd_pr__pfet_01v8__rdsw_diff_36 = 0.0
+ sky130_fd_pr__pfet_01v8__kt1_diff_36 = 0.0
+ sky130_fd_pr__pfet_01v8__pclm_diff_36 = 0.0
+ sky130_fd_pr__pfet_01v8__b0_diff_36 = -9.7759e-9
*
* sky130_fd_pr__pfet_01v8, Bin 037, W = 0.42, L = 2.0
* ----------------------------------
+ sky130_fd_pr__pfet_01v8__b0_diff_37 = -2.3998e-8
+ sky130_fd_pr__pfet_01v8__agidl_diff_37 = 0.0
+ sky130_fd_pr__pfet_01v8__b1_diff_37 = 6.7881e-9
+ sky130_fd_pr__pfet_01v8__ua_diff_37 = -7.2077e-12
+ sky130_fd_pr__pfet_01v8__bgidl_diff_37 = 0.0
+ sky130_fd_pr__pfet_01v8__nfactor_diff_37 = 0.4232
+ sky130_fd_pr__pfet_01v8__ub_diff_37 = 7.308e-19
+ sky130_fd_pr__pfet_01v8__tvoff_diff_37 = 0.0
+ sky130_fd_pr__pfet_01v8__ags_diff_37 = 0.0
+ sky130_fd_pr__pfet_01v8__k2_diff_37 = -0.0068908
+ sky130_fd_pr__pfet_01v8__pdits_diff_37 = 0.0
+ sky130_fd_pr__pfet_01v8__voff_diff_37 = -0.14578
+ sky130_fd_pr__pfet_01v8__eta0_diff_37 = 0.0
+ sky130_fd_pr__pfet_01v8__a0_diff_37 = 0.0
+ sky130_fd_pr__pfet_01v8__pditsd_diff_37 = 0.0
+ sky130_fd_pr__pfet_01v8__u0_diff_37 = 0.0032114
+ sky130_fd_pr__pfet_01v8__vsat_diff_37 = 0.0
+ sky130_fd_pr__pfet_01v8__vth0_diff_37 = 0.032454
+ sky130_fd_pr__pfet_01v8__cgidl_diff_37 = 0.0
+ sky130_fd_pr__pfet_01v8__keta_diff_37 = 0.0
+ sky130_fd_pr__pfet_01v8__rdsw_diff_37 = 0.0
+ sky130_fd_pr__pfet_01v8__kt1_diff_37 = 0.0
+ sky130_fd_pr__pfet_01v8__pclm_diff_37 = 0.0
*
* sky130_fd_pr__pfet_01v8, Bin 038, W = 0.42, L = 4.0
* ----------------------------------
+ sky130_fd_pr__pfet_01v8__pclm_diff_38 = 0.0
+ sky130_fd_pr__pfet_01v8__b0_diff_38 = -5.0871e-8
+ sky130_fd_pr__pfet_01v8__agidl_diff_38 = 0.0
+ sky130_fd_pr__pfet_01v8__b1_diff_38 = 1.1561e-9
+ sky130_fd_pr__pfet_01v8__ua_diff_38 = -3.8513e-13
+ sky130_fd_pr__pfet_01v8__bgidl_diff_38 = 0.0
+ sky130_fd_pr__pfet_01v8__nfactor_diff_38 = 0.46859
+ sky130_fd_pr__pfet_01v8__tvoff_diff_38 = 0.0
+ sky130_fd_pr__pfet_01v8__ags_diff_38 = 0.0
+ sky130_fd_pr__pfet_01v8__ub_diff_38 = 6.0269e-19
+ sky130_fd_pr__pfet_01v8__k2_diff_38 = -0.012379
+ sky130_fd_pr__pfet_01v8__pdits_diff_38 = 0.0
+ sky130_fd_pr__pfet_01v8__voff_diff_38 = -0.13346
+ sky130_fd_pr__pfet_01v8__eta0_diff_38 = 0.0
+ sky130_fd_pr__pfet_01v8__a0_diff_38 = 0.0
+ sky130_fd_pr__pfet_01v8__pditsd_diff_38 = 0.0
+ sky130_fd_pr__pfet_01v8__u0_diff_38 = 0.0029621
+ sky130_fd_pr__pfet_01v8__vsat_diff_38 = 0.0
+ sky130_fd_pr__pfet_01v8__vth0_diff_38 = 0.00040418
+ sky130_fd_pr__pfet_01v8__cgidl_diff_38 = 0.0
+ sky130_fd_pr__pfet_01v8__keta_diff_38 = 0.0
+ sky130_fd_pr__pfet_01v8__rdsw_diff_38 = 0.0
+ sky130_fd_pr__pfet_01v8__kt1_diff_38 = 0.0
*
* sky130_fd_pr__pfet_01v8, Bin 039, W = 0.42, L = 8.0
* ----------------------------------
+ sky130_fd_pr__pfet_01v8__kt1_diff_39 = 0.0
+ sky130_fd_pr__pfet_01v8__pclm_diff_39 = 0.0
+ sky130_fd_pr__pfet_01v8__b0_diff_39 = 1.4259e-7
+ sky130_fd_pr__pfet_01v8__agidl_diff_39 = 0.0
+ sky130_fd_pr__pfet_01v8__b1_diff_39 = -3.0094e-9
+ sky130_fd_pr__pfet_01v8__bgidl_diff_39 = 0.0
+ sky130_fd_pr__pfet_01v8__nfactor_diff_39 = 0.033193
+ sky130_fd_pr__pfet_01v8__ua_diff_39 = -1.1205e-11
+ sky130_fd_pr__pfet_01v8__tvoff_diff_39 = 0.0
+ sky130_fd_pr__pfet_01v8__ags_diff_39 = 0.0
+ sky130_fd_pr__pfet_01v8__ub_diff_39 = -2.7333e-20
+ sky130_fd_pr__pfet_01v8__k2_diff_39 = 0.0093948
+ sky130_fd_pr__pfet_01v8__pdits_diff_39 = 0.0
+ sky130_fd_pr__pfet_01v8__voff_diff_39 = -0.059118
+ sky130_fd_pr__pfet_01v8__eta0_diff_39 = 0.0
+ sky130_fd_pr__pfet_01v8__a0_diff_39 = 0.0
+ sky130_fd_pr__pfet_01v8__pditsd_diff_39 = 0.0
+ sky130_fd_pr__pfet_01v8__u0_diff_39 = -0.00034581
+ sky130_fd_pr__pfet_01v8__vsat_diff_39 = 0.0
+ sky130_fd_pr__pfet_01v8__vth0_diff_39 = 0.065303
+ sky130_fd_pr__pfet_01v8__cgidl_diff_39 = 0.0
+ sky130_fd_pr__pfet_01v8__keta_diff_39 = 0.0
+ sky130_fd_pr__pfet_01v8__rdsw_diff_39 = 0.0
*
* sky130_fd_pr__pfet_01v8, Bin 040, W = 0.42, L = 0.15
* -----------------------------------
+ sky130_fd_pr__pfet_01v8__rdsw_diff_40 = 0.0
+ sky130_fd_pr__pfet_01v8__kt1_diff_40 = 0.0
+ sky130_fd_pr__pfet_01v8__pclm_diff_40 = 0.0
+ sky130_fd_pr__pfet_01v8__b0_diff_40 = 3.2204e-7
+ sky130_fd_pr__pfet_01v8__b1_diff_40 = 2.0586e-8
+ sky130_fd_pr__pfet_01v8__agidl_diff_40 = 0.0
+ sky130_fd_pr__pfet_01v8__ua_diff_40 = -7.7662e-11
+ sky130_fd_pr__pfet_01v8__bgidl_diff_40 = 0.0
+ sky130_fd_pr__pfet_01v8__nfactor_diff_40 = 3.9999
+ sky130_fd_pr__pfet_01v8__ub_diff_40 = 6.1327e-19
+ sky130_fd_pr__pfet_01v8__pdits_diff_40 = 0.0
+ sky130_fd_pr__pfet_01v8__tvoff_diff_40 = 0.0
+ sky130_fd_pr__pfet_01v8__ags_diff_40 = 0.0
+ sky130_fd_pr__pfet_01v8__k2_diff_40 = -0.0067948
+ sky130_fd_pr__pfet_01v8__voff_diff_40 = -0.22293
+ sky130_fd_pr__pfet_01v8__a0_diff_40 = 0.0
+ sky130_fd_pr__pfet_01v8__pditsd_diff_40 = 0.0
+ sky130_fd_pr__pfet_01v8__eta0_diff_40 = 0.0
+ sky130_fd_pr__pfet_01v8__vsat_diff_40 = 18192.0
+ sky130_fd_pr__pfet_01v8__u0_diff_40 = 0.00058827
+ sky130_fd_pr__pfet_01v8__vth0_diff_40 = 0.010999
+ sky130_fd_pr__pfet_01v8__cgidl_diff_40 = 0.0
+ sky130_fd_pr__pfet_01v8__keta_diff_40 = 0.0
*
* sky130_fd_pr__pfet_01v8, Bin 041, W = 0.42, L = 0.18
* -----------------------------------
+ sky130_fd_pr__pfet_01v8__cgidl_diff_41 = 0.0
+ sky130_fd_pr__pfet_01v8__keta_diff_41 = 0.0
+ sky130_fd_pr__pfet_01v8__rdsw_diff_41 = 0.0
+ sky130_fd_pr__pfet_01v8__kt1_diff_41 = 0.0
+ sky130_fd_pr__pfet_01v8__pclm_diff_41 = 0.0
+ sky130_fd_pr__pfet_01v8__b0_diff_41 = -5.0000e-10
+ sky130_fd_pr__pfet_01v8__b1_diff_41 = 7.5436e-11
+ sky130_fd_pr__pfet_01v8__agidl_diff_41 = 0.0
+ sky130_fd_pr__pfet_01v8__ua_diff_41 = 8.8756e-10
+ sky130_fd_pr__pfet_01v8__bgidl_diff_41 = 0.0
+ sky130_fd_pr__pfet_01v8__nfactor_diff_41 = 5.1904
+ sky130_fd_pr__pfet_01v8__ub_diff_41 = 3.0505e-19
+ sky130_fd_pr__pfet_01v8__pdits_diff_41 = 0.0
+ sky130_fd_pr__pfet_01v8__tvoff_diff_41 = 0.0
+ sky130_fd_pr__pfet_01v8__ags_diff_41 = 0.0
+ sky130_fd_pr__pfet_01v8__k2_diff_41 = -2.5250e-2
+ sky130_fd_pr__pfet_01v8__voff_diff_41 = -0.25195
+ sky130_fd_pr__pfet_01v8__a0_diff_41 = 0.0
+ sky130_fd_pr__pfet_01v8__pditsd_diff_41 = 0.0
+ sky130_fd_pr__pfet_01v8__eta0_diff_41 = 0.0
+ sky130_fd_pr__pfet_01v8__vsat_diff_41 = 20962.0
+ sky130_fd_pr__pfet_01v8__u0_diff_41 = 4.2918e-3
+ sky130_fd_pr__pfet_01v8__vth0_diff_41 = -1.0000e-3
*
* sky130_fd_pr__pfet_01v8, Bin 042, W = 0.42, L = 0.5
* ----------------------------------
+ sky130_fd_pr__pfet_01v8__u0_diff_42 = 0.0018823
+ sky130_fd_pr__pfet_01v8__vth0_diff_42 = 0.037859
+ sky130_fd_pr__pfet_01v8__cgidl_diff_42 = 0.0
+ sky130_fd_pr__pfet_01v8__keta_diff_42 = 0.0
+ sky130_fd_pr__pfet_01v8__rdsw_diff_42 = 0.0
+ sky130_fd_pr__pfet_01v8__kt1_diff_42 = 0.0
+ sky130_fd_pr__pfet_01v8__pclm_diff_42 = 0.0
+ sky130_fd_pr__pfet_01v8__b0_diff_42 = 3.6809e-8
+ sky130_fd_pr__pfet_01v8__b1_diff_42 = -2.2779e-9
+ sky130_fd_pr__pfet_01v8__agidl_diff_42 = 0.0
+ sky130_fd_pr__pfet_01v8__ua_diff_42 = -1.0153e-11
+ sky130_fd_pr__pfet_01v8__bgidl_diff_42 = 0.0
+ sky130_fd_pr__pfet_01v8__nfactor_diff_42 = 0.98646
+ sky130_fd_pr__pfet_01v8__ub_diff_42 = 5.6326e-19
+ sky130_fd_pr__pfet_01v8__pdits_diff_42 = 0.0
+ sky130_fd_pr__pfet_01v8__tvoff_diff_42 = 0.0
+ sky130_fd_pr__pfet_01v8__ags_diff_42 = 0.0
+ sky130_fd_pr__pfet_01v8__k2_diff_42 = -0.0070988
+ sky130_fd_pr__pfet_01v8__voff_diff_42 = -0.21141
+ sky130_fd_pr__pfet_01v8__a0_diff_42 = 0.0
+ sky130_fd_pr__pfet_01v8__pditsd_diff_42 = 0.0
+ sky130_fd_pr__pfet_01v8__eta0_diff_42 = 0.0
+ sky130_fd_pr__pfet_01v8__vsat_diff_42 = 19837.0
*
* sky130_fd_pr__pfet_01v8, Bin 043, W = 0.55, L = 1.0
* ----------------------------------
+ sky130_fd_pr__pfet_01v8__pditsd_diff_43 = 0.0
+ sky130_fd_pr__pfet_01v8__eta0_diff_43 = 0.0
+ sky130_fd_pr__pfet_01v8__vsat_diff_43 = 119930.0
+ sky130_fd_pr__pfet_01v8__u0_diff_43 = 4.4042e-3
+ sky130_fd_pr__pfet_01v8__vth0_diff_43 = -1.1170e-2
+ sky130_fd_pr__pfet_01v8__cgidl_diff_43 = 0.0
+ sky130_fd_pr__pfet_01v8__keta_diff_43 = 0.0
+ sky130_fd_pr__pfet_01v8__rdsw_diff_43 = 0.0
+ sky130_fd_pr__pfet_01v8__kt1_diff_43 = 0.0
+ sky130_fd_pr__pfet_01v8__pclm_diff_43 = 0.0
+ sky130_fd_pr__pfet_01v8__b0_diff_43 = 1.2359e-7
+ sky130_fd_pr__pfet_01v8__b1_diff_43 = -2.1191e-9
+ sky130_fd_pr__pfet_01v8__agidl_diff_43 = 0.0
+ sky130_fd_pr__pfet_01v8__ua_diff_43 = 6.3881e-10
+ sky130_fd_pr__pfet_01v8__bgidl_diff_43 = 0.0
+ sky130_fd_pr__pfet_01v8__nfactor_diff_43 = 3.3479
+ sky130_fd_pr__pfet_01v8__ub_diff_43 = 6.1280e-21
+ sky130_fd_pr__pfet_01v8__pdits_diff_43 = 0.0
+ sky130_fd_pr__pfet_01v8__tvoff_diff_43 = 0.0
+ sky130_fd_pr__pfet_01v8__ags_diff_43 = 0.0
+ sky130_fd_pr__pfet_01v8__k2_diff_43 = -1.5500e-2
+ sky130_fd_pr__pfet_01v8__voff_diff_43 = -0.076218
+ sky130_fd_pr__pfet_01v8__a0_diff_43 = 0.0
*
* sky130_fd_pr__pfet_01v8, Bin 044, W = 0.55, L = 2.0
* ----------------------------------
+ sky130_fd_pr__pfet_01v8__voff_diff_44 = -0.11697
+ sky130_fd_pr__pfet_01v8__a0_diff_44 = 0.0
+ sky130_fd_pr__pfet_01v8__pditsd_diff_44 = 0.0
+ sky130_fd_pr__pfet_01v8__eta0_diff_44 = 0.0
+ sky130_fd_pr__pfet_01v8__vsat_diff_44 = 0.0
+ sky130_fd_pr__pfet_01v8__u0_diff_44 = 0.0030762
+ sky130_fd_pr__pfet_01v8__vth0_diff_44 = 0.027087
+ sky130_fd_pr__pfet_01v8__cgidl_diff_44 = 0.0
+ sky130_fd_pr__pfet_01v8__keta_diff_44 = 0.0
+ sky130_fd_pr__pfet_01v8__rdsw_diff_44 = 0.0
+ sky130_fd_pr__pfet_01v8__kt1_diff_44 = 0.0
+ sky130_fd_pr__pfet_01v8__pclm_diff_44 = 0.0
+ sky130_fd_pr__pfet_01v8__b0_diff_44 = -1.9488e-8
+ sky130_fd_pr__pfet_01v8__b1_diff_44 = 3.5905e-10
+ sky130_fd_pr__pfet_01v8__agidl_diff_44 = 0.0
+ sky130_fd_pr__pfet_01v8__ua_diff_44 = 9.5215e-12
+ sky130_fd_pr__pfet_01v8__bgidl_diff_44 = 0.0
+ sky130_fd_pr__pfet_01v8__nfactor_diff_44 = 0.31697
+ sky130_fd_pr__pfet_01v8__ub_diff_44 = 6.6875e-19
+ sky130_fd_pr__pfet_01v8__pdits_diff_44 = 0.0
+ sky130_fd_pr__pfet_01v8__tvoff_diff_44 = 0.0
+ sky130_fd_pr__pfet_01v8__ags_diff_44 = 0.0
+ sky130_fd_pr__pfet_01v8__k2_diff_44 = -0.0090663
*
* sky130_fd_pr__pfet_01v8, Bin 045, W = 0.55, L = 4.0
* ----------------------------------
+ sky130_fd_pr__pfet_01v8__pdits_diff_45 = 0.0
+ sky130_fd_pr__pfet_01v8__tvoff_diff_45 = 0.0
+ sky130_fd_pr__pfet_01v8__ags_diff_45 = 0.0
+ sky130_fd_pr__pfet_01v8__k2_diff_45 = 0.01045
+ sky130_fd_pr__pfet_01v8__voff_diff_45 = -0.059301
+ sky130_fd_pr__pfet_01v8__a0_diff_45 = 0.0
+ sky130_fd_pr__pfet_01v8__pditsd_diff_45 = 0.0
+ sky130_fd_pr__pfet_01v8__eta0_diff_45 = 0.0
+ sky130_fd_pr__pfet_01v8__vsat_diff_45 = 0.0
+ sky130_fd_pr__pfet_01v8__u0_diff_45 = -0.00056442
+ sky130_fd_pr__pfet_01v8__vth0_diff_45 = 0.067926
+ sky130_fd_pr__pfet_01v8__cgidl_diff_45 = 0.0
+ sky130_fd_pr__pfet_01v8__keta_diff_45 = 0.0
+ sky130_fd_pr__pfet_01v8__rdsw_diff_45 = 0.0
+ sky130_fd_pr__pfet_01v8__kt1_diff_45 = 0.0
+ sky130_fd_pr__pfet_01v8__pclm_diff_45 = 0.0
+ sky130_fd_pr__pfet_01v8__b0_diff_45 = 9.2682e-8
+ sky130_fd_pr__pfet_01v8__b1_diff_45 = -3.0393e-10
+ sky130_fd_pr__pfet_01v8__agidl_diff_45 = 0.0
+ sky130_fd_pr__pfet_01v8__ua_diff_45 = -9.3232e-12
+ sky130_fd_pr__pfet_01v8__bgidl_diff_45 = 0.0
+ sky130_fd_pr__pfet_01v8__nfactor_diff_45 = -0.21757
+ sky130_fd_pr__pfet_01v8__ub_diff_45 = -3.8525e-20
*
* sky130_fd_pr__pfet_01v8, Bin 046, W = 0.55, L = 8.0
* ----------------------------------
+ sky130_fd_pr__pfet_01v8__bgidl_diff_46 = 0.0
+ sky130_fd_pr__pfet_01v8__nfactor_diff_46 = 0.59995
+ sky130_fd_pr__pfet_01v8__ub_diff_46 = 6.9222e-19
+ sky130_fd_pr__pfet_01v8__pdits_diff_46 = 0.0
+ sky130_fd_pr__pfet_01v8__tvoff_diff_46 = 0.0
+ sky130_fd_pr__pfet_01v8__ags_diff_46 = 0.0
+ sky130_fd_pr__pfet_01v8__k2_diff_46 = -0.013366
+ sky130_fd_pr__pfet_01v8__voff_diff_46 = -0.14278
+ sky130_fd_pr__pfet_01v8__a0_diff_46 = 0.0
+ sky130_fd_pr__pfet_01v8__eta0_diff_46 = 0.0
+ sky130_fd_pr__pfet_01v8__pditsd_diff_46 = 0.0
+ sky130_fd_pr__pfet_01v8__u0_diff_46 = 0.0034898
+ sky130_fd_pr__pfet_01v8__vsat_diff_46 = 0.0
+ sky130_fd_pr__pfet_01v8__vth0_diff_46 = 0.0039578
+ sky130_fd_pr__pfet_01v8__cgidl_diff_46 = 0.0
+ sky130_fd_pr__pfet_01v8__keta_diff_46 = 0.0
+ sky130_fd_pr__pfet_01v8__rdsw_diff_46 = 0.0
+ sky130_fd_pr__pfet_01v8__kt1_diff_46 = 0.0
+ sky130_fd_pr__pfet_01v8__pclm_diff_46 = 0.0
+ sky130_fd_pr__pfet_01v8__b0_diff_46 = -2.1309e-8
+ sky130_fd_pr__pfet_01v8__b1_diff_46 = 2.2477e-9
+ sky130_fd_pr__pfet_01v8__agidl_diff_46 = 0.0
+ sky130_fd_pr__pfet_01v8__ua_diff_46 = -2.4775e-12
*
* sky130_fd_pr__pfet_01v8, Bin 047, W = 0.55, L = 0.15
* -----------------------------------
+ sky130_fd_pr__pfet_01v8__agidl_diff_47 = 0.0
+ sky130_fd_pr__pfet_01v8__b1_diff_47 = 2.3324e-8
+ sky130_fd_pr__pfet_01v8__ua_diff_47 = -4.2037e-11
+ sky130_fd_pr__pfet_01v8__bgidl_diff_47 = 0.0
+ sky130_fd_pr__pfet_01v8__nfactor_diff_47 = 3.9781
+ sky130_fd_pr__pfet_01v8__ub_diff_47 = 5.792e-19
+ sky130_fd_pr__pfet_01v8__pdits_diff_47 = 0.0
+ sky130_fd_pr__pfet_01v8__tvoff_diff_47 = 0.0
+ sky130_fd_pr__pfet_01v8__ags_diff_47 = 0.0
+ sky130_fd_pr__pfet_01v8__k2_diff_47 = 0.0089906
+ sky130_fd_pr__pfet_01v8__voff_diff_47 = -0.22208
+ sky130_fd_pr__pfet_01v8__eta0_diff_47 = 0.0
+ sky130_fd_pr__pfet_01v8__a0_diff_47 = 0.0
+ sky130_fd_pr__pfet_01v8__pditsd_diff_47 = 0.0
+ sky130_fd_pr__pfet_01v8__u0_diff_47 = 0.00068298
+ sky130_fd_pr__pfet_01v8__vsat_diff_47 = 21559.0
+ sky130_fd_pr__pfet_01v8__vth0_diff_47 = -0.013366
+ sky130_fd_pr__pfet_01v8__cgidl_diff_47 = 0.0
+ sky130_fd_pr__pfet_01v8__keta_diff_47 = 0.0
+ sky130_fd_pr__pfet_01v8__rdsw_diff_47 = 0.0
+ sky130_fd_pr__pfet_01v8__kt1_diff_47 = 0.0
+ sky130_fd_pr__pfet_01v8__pclm_diff_47 = 0.0
+ sky130_fd_pr__pfet_01v8__b0_diff_47 = 6.8027e-7
*
* sky130_fd_pr__pfet_01v8, Bin 048, W = 0.55, L = 0.5
* ----------------------------------
+ sky130_fd_pr__pfet_01v8__b0_diff_48 = 2.4391e-8
+ sky130_fd_pr__pfet_01v8__agidl_diff_48 = 0.0
+ sky130_fd_pr__pfet_01v8__b1_diff_48 = 1.6514e-8
+ sky130_fd_pr__pfet_01v8__ua_diff_48 = -4.9634e-12
+ sky130_fd_pr__pfet_01v8__bgidl_diff_48 = 0.0
+ sky130_fd_pr__pfet_01v8__nfactor_diff_48 = 0.48298
+ sky130_fd_pr__pfet_01v8__ub_diff_48 = 4.8904e-19
+ sky130_fd_pr__pfet_01v8__tvoff_diff_48 = 0.0
+ sky130_fd_pr__pfet_01v8__ags_diff_48 = 0.0
+ sky130_fd_pr__pfet_01v8__k2_diff_48 = -0.016336
+ sky130_fd_pr__pfet_01v8__pdits_diff_48 = 0.0
+ sky130_fd_pr__pfet_01v8__voff_diff_48 = -0.17412
+ sky130_fd_pr__pfet_01v8__eta0_diff_48 = 0.0
+ sky130_fd_pr__pfet_01v8__a0_diff_48 = 0.0
+ sky130_fd_pr__pfet_01v8__pditsd_diff_48 = 0.0
+ sky130_fd_pr__pfet_01v8__u0_diff_48 = 0.0015741
+ sky130_fd_pr__pfet_01v8__vsat_diff_48 = 19810.0
+ sky130_fd_pr__pfet_01v8__vth0_diff_48 = 0.038899
+ sky130_fd_pr__pfet_01v8__cgidl_diff_48 = 0.0
+ sky130_fd_pr__pfet_01v8__keta_diff_48 = 0.0
+ sky130_fd_pr__pfet_01v8__rdsw_diff_48 = 0.0
+ sky130_fd_pr__pfet_01v8__kt1_diff_48 = 0.0
+ sky130_fd_pr__pfet_01v8__pclm_diff_48 = 0.0
*
* sky130_fd_pr__pfet_01v8, Bin 049, W = 0.64, L = 0.15
* -----------------------------------
+ sky130_fd_pr__pfet_01v8__pclm_diff_49 = 0.0
+ sky130_fd_pr__pfet_01v8__b0_diff_49 = 8.6951e-7
+ sky130_fd_pr__pfet_01v8__agidl_diff_49 = 0.0
+ sky130_fd_pr__pfet_01v8__b1_diff_49 = 9.8831e-9
+ sky130_fd_pr__pfet_01v8__ua_diff_49 = -2.0555e-10
+ sky130_fd_pr__pfet_01v8__bgidl_diff_49 = 0.0
+ sky130_fd_pr__pfet_01v8__nfactor_diff_49 = 4.0
+ sky130_fd_pr__pfet_01v8__tvoff_diff_49 = 0.0
+ sky130_fd_pr__pfet_01v8__ags_diff_49 = 0.0
+ sky130_fd_pr__pfet_01v8__ub_diff_49 = 6.2299e-19
+ sky130_fd_pr__pfet_01v8__k2_diff_49 = 0.014274
+ sky130_fd_pr__pfet_01v8__pdits_diff_49 = 0.0
+ sky130_fd_pr__pfet_01v8__voff_diff_49 = -0.17738
+ sky130_fd_pr__pfet_01v8__eta0_diff_49 = 0.0
+ sky130_fd_pr__pfet_01v8__a0_diff_49 = 0.0
+ sky130_fd_pr__pfet_01v8__pditsd_diff_49 = 0.0
+ sky130_fd_pr__pfet_01v8__u0_diff_49 = 0.0001875
+ sky130_fd_pr__pfet_01v8__vsat_diff_49 = 24231.0
+ sky130_fd_pr__pfet_01v8__vth0_diff_49 = -0.10266
+ sky130_fd_pr__pfet_01v8__cgidl_diff_49 = 0.0
+ sky130_fd_pr__pfet_01v8__keta_diff_49 = 0.0
+ sky130_fd_pr__pfet_01v8__rdsw_diff_49 = 0.0
+ sky130_fd_pr__pfet_01v8__kt1_diff_49 = 0.0
*
* sky130_fd_pr__pfet_01v8, Bin 050, W = 0.84, L = 0.15
* -----------------------------------
+ sky130_fd_pr__pfet_01v8__kt1_diff_50 = 0.0
+ sky130_fd_pr__pfet_01v8__pclm_diff_50 = 0.0
+ sky130_fd_pr__pfet_01v8__b0_diff_50 = 0.0
+ sky130_fd_pr__pfet_01v8__b1_diff_50 = 0.0
+ sky130_fd_pr__pfet_01v8__agidl_diff_50 = 0.0
+ sky130_fd_pr__pfet_01v8__ua_diff_50 = -2.4122e-10
+ sky130_fd_pr__pfet_01v8__bgidl_diff_50 = 0.0
+ sky130_fd_pr__pfet_01v8__nfactor_diff_50 = 3.5042
+ sky130_fd_pr__pfet_01v8__ub_diff_50 = 6.4451e-19
+ sky130_fd_pr__pfet_01v8__pdits_diff_50 = 0.0
+ sky130_fd_pr__pfet_01v8__tvoff_diff_50 = 0.0
+ sky130_fd_pr__pfet_01v8__ags_diff_50 = 0.0
+ sky130_fd_pr__pfet_01v8__k2_diff_50 = -0.024696
+ sky130_fd_pr__pfet_01v8__voff_diff_50 = -0.15812
+ sky130_fd_pr__pfet_01v8__a0_diff_50 = 0.0
+ sky130_fd_pr__pfet_01v8__pditsd_diff_50 = 0.0
+ sky130_fd_pr__pfet_01v8__eta0_diff_50 = 0.0
+ sky130_fd_pr__pfet_01v8__vsat_diff_50 = -20000.0
+ sky130_fd_pr__pfet_01v8__u0_diff_50 = 0.00027636
+ sky130_fd_pr__pfet_01v8__vth0_diff_50 = -0.12447
+ sky130_fd_pr__pfet_01v8__cgidl_diff_50 = 0.0
+ sky130_fd_pr__pfet_01v8__keta_diff_50 = 0.0
+ sky130_fd_pr__pfet_01v8__rdsw_diff_50 = 0.0
*
* sky130_fd_pr__pfet_01v8, Bin 051, W = 1.65, L = 0.15
* -----------------------------------
+ sky130_fd_pr__pfet_01v8__rdsw_diff_51 = 0.0
+ sky130_fd_pr__pfet_01v8__kt1_diff_51 = 0.0
+ sky130_fd_pr__pfet_01v8__pclm_diff_51 = 0.0
+ sky130_fd_pr__pfet_01v8__b0_diff_51 = 0.0
+ sky130_fd_pr__pfet_01v8__b1_diff_51 = 0.0
+ sky130_fd_pr__pfet_01v8__agidl_diff_51 = 0.0
+ sky130_fd_pr__pfet_01v8__ua_diff_51 = -2.8822e-11
+ sky130_fd_pr__pfet_01v8__bgidl_diff_51 = 0.0
+ sky130_fd_pr__pfet_01v8__nfactor_diff_51 = 2.8705
+ sky130_fd_pr__pfet_01v8__ub_diff_51 = 3.1525e-19
+ sky130_fd_pr__pfet_01v8__pdits_diff_51 = 0.0
+ sky130_fd_pr__pfet_01v8__tvoff_diff_51 = 0.0
+ sky130_fd_pr__pfet_01v8__ags_diff_51 = 0.0
+ sky130_fd_pr__pfet_01v8__k2_diff_51 = -0.0044952
+ sky130_fd_pr__pfet_01v8__voff_diff_51 = -0.21797
+ sky130_fd_pr__pfet_01v8__a0_diff_51 = 0.0
+ sky130_fd_pr__pfet_01v8__pditsd_diff_51 = 0.0
+ sky130_fd_pr__pfet_01v8__eta0_diff_51 = 0.0
+ sky130_fd_pr__pfet_01v8__vsat_diff_51 = -16774.0
+ sky130_fd_pr__pfet_01v8__u0_diff_51 = 0.00036783
+ sky130_fd_pr__pfet_01v8__vth0_diff_51 = -0.10906
+ sky130_fd_pr__pfet_01v8__cgidl_diff_51 = 0.0
+ sky130_fd_pr__pfet_01v8__keta_diff_51 = 0.0
.include "sky130_fd_pr__pfet_01v8.pm3.spice"
