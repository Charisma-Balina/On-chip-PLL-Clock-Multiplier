* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.

* SKY130 Spice File.
.param
+ sky130_fd_pr__nfet_20v0__nwgatejunction_mult=7.5058e-01
+ sky130_fd_pr__nfet_20v0__nwgatemjswjunction_mult = 8.3390e-1
+ sky130_fd_pr__nfet_20v0__nwgatepbswjunction_mult = 1.0204e+0
+ sky130_fd_pr__nfet_20v0__nwgatectjunction_mult = 1.0
+ sky130_fd_pr__nfet_20v0_iso__vb = 26.0
.model sky130_fd_pr__model__parasitic__diode_pw2dn__extended_drain d
+ level = 3.0
+ tlevc = 1.0
+ scalm = 1.0e-6
+ area = 1.0e+12
* Junction Capacitance Parameters
+ cj = '0.00038945*sky130_fd_pr__nfet_20v0__nwgatejunction_mult*1e-12*sky130_fd_pr__model__parasitic__diode_pw2dn__ajunction_mult' $ Units: farad/meter^2
+ mj = '0.63982*sky130_fd_pr__nfet_20v0__nwgatemjswjunction_mult'
+ pb = '0.58758*sky130_fd_pr__nfet_20v0__nwgatepbswjunction_mult' $ Units: volt
+ cjsw = '3.743e-010*sky130_fd_pr__nfet_20v0__nwgatejunction_mult*1e-6*sky130_fd_pr__model__parasitic__diode_pw2dn__pjunction_mult' $ Units: farad/meter
+ mjsw = '0.80357*sky130_fd_pr__nfet_20v0__nwgatemjswjunction_mult'
+ php = '0.2500*sky130_fd_pr__nfet_20v0__nwgatepbswjunction_mult' $ Units: volt
+ cta = '0.0016157*sky130_fd_pr__nfet_20v0__nwgatectjunction_mult' $ Units: 1/coulomb
+ ctp = '0.0008*sky130_fd_pr__nfet_20v0__nwgatectjunction_mult' $ Units: 1/coulomb
+ tpb = 0.0010003 $ Units: volt/coulomb
+ tphp = 0.000675 $ Units: volt/coulomb
* Diode IV Parameters
+ js = 1.4693e-017 $ Units: amper/meter^2
+ jsw = 7.41e-018 $ Units: amper/meter
+ n = 1.0791
+ rs = 900 $ Units: ohm (ohm/meter^2 if area defined)
+ ik = '2.08e-009/1e-12' $ Units: amper/meter^2
+ ikr = '0/1e-12' $ Units: amper/meter^2
+ vb = 'sky130_fd_pr__nfet_20v0_iso__vb' $ Units: volt
+ ibv = 0.00106 $ Units: amper
+ trs = 0 $ Units: 1/coulomb
+ xti = 3.0
+ eg = 1.50 $ Units: electron-volt
+ tref = 30 $ Units: coulomb
* Default Parameters
+ tcv = 0 $ Units: 1/coulomb
+ gap1 = 0.000473 $ Units: electron-volt/coulomb
+ gap2 = 1110.0
+ ttt1 = 0 $ Units: 1/coulomb
+ ttt2 = 0 $ Units: 1/coulomb^2
+ tm1 = 0 $ Units: 1/coulomb
+ tm2 = 0 $ Units: 1/coulomb^2
+ lm = 0 $ Units: meter
+ lp = 0 $ Units: meter
+ wm = 0 $ Units: meter
+ wp = 0 $ Units: meter
+ xm = 0 $ Units: meter
+ xoi = 10000.0
+ xom = 10000 $ Units: angstrom
+ xp = 0 $ Units: meter
+ xw = 0 $ Units: meter
