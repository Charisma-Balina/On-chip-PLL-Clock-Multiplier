magic
tech sky130A
timestamp 1605977318
<< nwell >>
rect 89 535 767 640
rect 137 479 767 535
rect 505 460 767 479
rect 677 307 767 308
rect 443 295 767 307
rect 397 157 767 295
rect 397 31 514 157
<< nmos >>
rect 70 397 310 412
rect 554 368 569 404
rect 70 341 250 356
rect 605 356 620 404
rect 70 284 106 299
rect 199 92 214 128
rect 256 92 271 272
rect 312 92 327 332
rect 579 83 594 119
rect 630 71 645 119
<< pmos >>
rect 155 530 220 545
rect 287 530 352 545
rect 554 502 569 574
rect 605 478 620 574
rect 448 207 463 272
rect 579 217 594 289
rect 630 193 645 289
rect 448 75 463 140
<< ndiff >>
rect 70 437 310 445
rect 70 420 99 437
rect 116 420 133 437
rect 150 420 167 437
rect 184 420 201 437
rect 218 420 235 437
rect 252 420 269 437
rect 286 420 310 437
rect 70 412 310 420
rect 70 389 310 397
rect 523 394 554 404
rect 70 372 74 389
rect 91 372 108 389
rect 125 372 142 389
rect 159 372 176 389
rect 193 372 210 389
rect 227 372 261 389
rect 278 372 310 389
rect 70 365 310 372
rect 523 377 529 394
rect 546 377 554 394
rect 523 368 554 377
rect 569 380 605 404
rect 569 368 582 380
rect 70 356 250 365
rect 70 308 250 341
rect 578 363 582 368
rect 599 363 605 380
rect 578 356 605 363
rect 620 389 649 404
rect 620 372 628 389
rect 645 372 649 389
rect 620 356 649 372
rect 280 317 312 332
rect 70 299 106 308
rect 280 300 287 317
rect 304 300 312 317
rect 70 276 106 284
rect 70 259 80 276
rect 97 259 106 276
rect 70 251 106 259
rect 280 283 312 300
rect 280 272 287 283
rect 223 128 256 272
rect 166 118 199 128
rect 166 101 174 118
rect 191 101 199 118
rect 166 92 199 101
rect 214 92 256 128
rect 271 266 287 272
rect 304 266 312 283
rect 271 249 312 266
rect 271 232 287 249
rect 304 232 312 249
rect 271 215 312 232
rect 271 198 287 215
rect 304 198 312 215
rect 271 181 312 198
rect 271 164 287 181
rect 304 164 312 181
rect 271 147 312 164
rect 271 130 287 147
rect 304 130 312 147
rect 271 113 312 130
rect 271 96 287 113
rect 304 96 312 113
rect 271 92 312 96
rect 327 301 360 332
rect 327 284 335 301
rect 352 284 360 301
rect 327 267 360 284
rect 327 250 335 267
rect 352 250 360 267
rect 327 215 360 250
rect 327 198 335 215
rect 352 198 360 215
rect 327 181 360 198
rect 327 164 335 181
rect 352 164 360 181
rect 327 147 360 164
rect 327 130 335 147
rect 352 130 360 147
rect 327 113 360 130
rect 327 96 335 113
rect 352 96 360 113
rect 327 92 360 96
rect 548 109 579 119
rect 548 92 554 109
rect 571 92 579 109
rect 548 83 579 92
rect 594 95 630 119
rect 594 83 607 95
rect 603 78 607 83
rect 624 78 630 95
rect 603 71 630 78
rect 645 104 674 119
rect 645 87 653 104
rect 670 87 674 104
rect 645 71 674 87
<< pdiff >>
rect 155 570 220 578
rect 155 553 159 570
rect 176 553 193 570
rect 210 553 220 570
rect 287 570 352 578
rect 155 545 220 553
rect 155 522 220 530
rect 155 505 163 522
rect 180 505 199 522
rect 216 505 220 522
rect 287 553 291 570
rect 308 553 325 570
rect 342 553 352 570
rect 287 545 352 553
rect 523 570 554 574
rect 523 553 529 570
rect 546 553 554 570
rect 523 536 554 553
rect 287 522 352 530
rect 155 497 220 505
rect 287 505 296 522
rect 313 505 330 522
rect 347 505 352 522
rect 287 497 352 505
rect 523 519 529 536
rect 546 519 554 536
rect 523 502 554 519
rect 569 570 605 574
rect 569 553 582 570
rect 599 553 605 570
rect 569 536 605 553
rect 569 519 582 536
rect 599 519 605 536
rect 569 502 605 519
rect 578 478 605 502
rect 620 570 650 574
rect 620 553 627 570
rect 644 553 650 570
rect 620 536 650 553
rect 620 519 627 536
rect 644 519 650 536
rect 620 478 650 519
rect 548 285 579 289
rect 415 267 448 272
rect 415 250 423 267
rect 440 250 448 267
rect 415 233 448 250
rect 415 216 423 233
rect 440 216 448 233
rect 415 207 448 216
rect 463 262 496 272
rect 463 245 471 262
rect 488 245 496 262
rect 463 228 496 245
rect 463 211 471 228
rect 488 211 496 228
rect 548 268 554 285
rect 571 268 579 285
rect 548 251 579 268
rect 548 234 554 251
rect 571 234 579 251
rect 548 217 579 234
rect 594 285 630 289
rect 594 268 607 285
rect 624 268 630 285
rect 594 251 630 268
rect 594 234 607 251
rect 624 234 630 251
rect 594 217 630 234
rect 463 207 496 211
rect 603 193 630 217
rect 645 285 675 289
rect 645 268 652 285
rect 669 268 675 285
rect 645 251 675 268
rect 645 234 652 251
rect 669 234 675 251
rect 645 193 675 234
rect 415 136 448 140
rect 415 119 423 136
rect 440 119 448 136
rect 415 100 448 119
rect 415 83 423 100
rect 440 83 448 100
rect 415 75 448 83
rect 463 130 496 140
rect 463 113 471 130
rect 488 113 496 130
rect 463 96 496 113
rect 463 79 471 96
rect 488 79 496 96
rect 463 75 496 79
<< ndiffc >>
rect 99 420 116 437
rect 133 420 150 437
rect 167 420 184 437
rect 201 420 218 437
rect 235 420 252 437
rect 269 420 286 437
rect 74 372 91 389
rect 108 372 125 389
rect 142 372 159 389
rect 176 372 193 389
rect 210 372 227 389
rect 261 372 278 389
rect 529 377 546 394
rect 582 363 599 380
rect 628 372 645 389
rect 287 300 304 317
rect 80 259 97 276
rect 174 101 191 118
rect 287 266 304 283
rect 287 232 304 249
rect 287 198 304 215
rect 287 164 304 181
rect 287 130 304 147
rect 287 96 304 113
rect 335 284 352 301
rect 335 250 352 267
rect 335 198 352 215
rect 335 164 352 181
rect 335 130 352 147
rect 335 96 352 113
rect 554 92 571 109
rect 607 78 624 95
rect 653 87 670 104
<< pdiffc >>
rect 159 553 176 570
rect 193 553 210 570
rect 163 505 180 522
rect 199 505 216 522
rect 291 553 308 570
rect 325 553 342 570
rect 529 553 546 570
rect 296 505 313 522
rect 330 505 347 522
rect 529 519 546 536
rect 582 553 599 570
rect 582 519 599 536
rect 627 553 644 570
rect 627 519 644 536
rect 423 250 440 267
rect 423 216 440 233
rect 471 245 488 262
rect 471 211 488 228
rect 554 268 571 285
rect 554 234 571 251
rect 607 268 624 285
rect 607 234 624 251
rect 652 268 669 285
rect 652 234 669 251
rect 423 119 440 136
rect 423 83 440 100
rect 471 113 488 130
rect 471 79 488 96
<< psubdiff >>
rect 448 393 460 410
rect 477 393 489 410
rect 448 392 489 393
rect 448 348 460 365
rect 477 348 489 365
rect 448 347 489 348
<< nsubdiff >>
rect 116 605 128 622
rect 145 605 157 622
rect 198 605 210 622
rect 227 605 239 622
rect 280 605 292 622
rect 309 605 321 622
rect 362 605 374 622
rect 391 605 403 622
rect 444 605 456 622
rect 473 605 485 622
rect 704 266 716 283
rect 733 266 745 283
rect 704 220 716 237
rect 733 220 745 237
rect 704 176 716 193
rect 733 176 745 193
<< psubdiffcont >>
rect 460 393 477 410
rect 460 348 477 365
<< nsubdiffcont >>
rect 128 605 145 622
rect 210 605 227 622
rect 292 605 309 622
rect 374 605 391 622
rect 456 605 473 622
rect 716 266 733 283
rect 716 220 733 237
rect 716 176 733 193
<< poly >>
rect 554 574 569 587
rect 605 574 620 587
rect 240 546 267 554
rect 240 545 245 546
rect 142 530 155 545
rect 220 530 245 545
rect 240 529 245 530
rect 262 545 267 546
rect 262 530 287 545
rect 352 530 365 545
rect 262 529 267 530
rect 240 521 267 529
rect 245 474 262 521
rect 245 459 340 474
rect 554 462 569 502
rect 605 468 620 478
rect 323 412 340 459
rect 541 457 569 462
rect 602 461 620 468
rect 538 440 546 457
rect 563 440 570 457
rect 591 452 620 461
rect 541 435 569 440
rect 46 397 70 412
rect 310 397 340 412
rect 46 356 61 397
rect 554 404 569 435
rect 591 435 596 452
rect 613 435 620 452
rect 591 427 620 435
rect 602 421 620 427
rect 605 404 620 421
rect 8 343 70 356
rect 8 326 13 343
rect 30 341 70 343
rect 250 341 263 356
rect 30 326 35 341
rect 8 318 35 326
rect 312 340 394 356
rect 554 353 569 368
rect 605 343 620 356
rect 312 332 327 340
rect 57 284 70 299
rect 106 284 271 299
rect 117 281 271 284
rect 117 228 132 281
rect 256 272 271 281
rect 90 223 132 228
rect 90 206 98 223
rect 115 206 132 223
rect 90 201 132 206
rect 176 168 214 173
rect 176 151 184 168
rect 201 151 214 168
rect 176 146 214 151
rect 199 128 214 146
rect 374 182 394 340
rect 579 289 594 302
rect 630 289 645 302
rect 448 272 463 285
rect 448 187 463 207
rect 439 182 472 187
rect 374 165 447 182
rect 464 165 472 182
rect 579 177 594 217
rect 630 183 645 193
rect 566 172 594 177
rect 627 176 645 183
rect 439 160 472 165
rect 448 140 463 160
rect 563 155 571 172
rect 588 155 595 172
rect 616 167 645 176
rect 566 150 594 155
rect 199 77 214 92
rect 256 83 271 92
rect 312 83 327 92
rect 256 68 327 83
rect 579 119 594 150
rect 616 150 621 167
rect 638 150 645 167
rect 616 142 645 150
rect 627 136 645 142
rect 630 119 645 136
rect 448 62 463 75
rect 579 68 594 83
rect 630 58 645 71
<< polycont >>
rect 245 529 262 546
rect 546 440 563 457
rect 596 435 613 452
rect 13 326 30 343
rect 98 206 115 223
rect 184 151 201 168
rect 447 165 464 182
rect 571 155 588 172
rect 621 150 638 167
<< locali >>
rect 0 605 80 622
rect 97 605 114 622
rect 145 605 148 622
rect 165 605 182 622
rect 199 605 210 622
rect 233 605 250 622
rect 267 605 284 622
rect 309 605 318 622
rect 335 605 352 622
rect 369 605 374 622
rect 403 605 420 622
rect 437 605 454 622
rect 473 605 488 622
rect 505 605 522 622
rect 539 605 556 622
rect 573 605 590 622
rect 607 605 624 622
rect 641 605 658 622
rect 675 605 767 622
rect 165 572 207 605
rect 151 570 222 572
rect 151 553 159 570
rect 176 553 193 570
rect 210 553 222 570
rect 151 551 222 553
rect 242 570 352 571
rect 242 553 291 570
rect 308 553 325 570
rect 342 553 352 570
rect 242 552 352 553
rect 526 570 548 578
rect 526 553 529 570
rect 546 553 548 570
rect 242 546 265 552
rect 242 529 245 546
rect 262 529 265 546
rect 155 522 224 524
rect 155 505 163 522
rect 180 505 199 522
rect 216 505 224 522
rect 242 521 265 529
rect 526 536 548 553
rect 284 522 355 523
rect 155 488 224 505
rect 37 463 224 488
rect 284 505 296 522
rect 313 505 330 522
rect 347 505 355 522
rect 284 504 355 505
rect 526 519 529 536
rect 546 519 548 536
rect 37 395 64 463
rect 284 457 328 504
rect 526 491 548 519
rect 577 570 600 605
rect 577 553 582 570
rect 599 553 600 570
rect 577 536 600 553
rect 577 519 582 536
rect 599 519 600 536
rect 577 508 600 519
rect 627 570 656 578
rect 644 553 656 570
rect 627 536 656 553
rect 644 519 656 536
rect 526 474 610 491
rect 627 478 656 519
rect 590 461 610 474
rect 284 445 546 457
rect 87 440 546 445
rect 563 440 571 457
rect 590 452 613 461
rect 87 437 329 440
rect 87 420 99 437
rect 116 420 133 437
rect 150 420 167 437
rect 184 420 201 437
rect 218 420 235 437
rect 252 420 269 437
rect 286 420 329 437
rect 590 435 596 452
rect 590 427 613 435
rect 590 423 609 427
rect 87 419 329 420
rect 37 389 310 395
rect 37 372 74 389
rect 91 372 108 389
rect 125 372 142 389
rect 159 372 176 389
rect 193 372 210 389
rect 227 372 261 389
rect 278 372 310 389
rect 37 371 310 372
rect 434 393 460 410
rect 477 393 501 410
rect 434 365 501 393
rect 525 406 609 423
rect 525 394 547 406
rect 639 404 656 478
rect 525 377 529 394
rect 546 377 547 394
rect 626 389 656 404
rect 525 368 547 377
rect 578 380 600 388
rect 4 343 31 351
rect 4 326 13 343
rect 30 326 31 343
rect 434 348 460 365
rect 477 348 501 365
rect 4 174 31 326
rect 286 317 305 332
rect 286 300 287 317
rect 304 300 305 317
rect 286 283 305 300
rect 78 276 99 278
rect 70 259 80 276
rect 97 259 106 276
rect 286 266 287 283
rect 304 266 305 283
rect 78 251 99 259
rect 286 249 305 266
rect 286 232 287 249
rect 304 232 305 249
rect 90 206 98 223
rect 115 206 123 223
rect 286 215 305 232
rect 286 198 287 215
rect 304 198 305 215
rect 286 181 305 198
rect 4 168 210 174
rect 4 151 184 168
rect 201 151 210 168
rect 4 145 210 151
rect 286 164 287 181
rect 304 164 305 181
rect 286 147 305 164
rect 173 118 191 128
rect 173 101 174 118
rect 173 92 191 101
rect 286 124 287 147
rect 304 124 305 147
rect 286 113 305 124
rect 286 96 287 113
rect 304 96 305 113
rect 286 86 305 96
rect 334 301 353 332
rect 434 329 501 348
rect 578 363 582 380
rect 599 363 600 380
rect 578 336 600 363
rect 626 372 628 389
rect 645 372 656 389
rect 626 356 656 372
rect 556 329 623 336
rect 434 312 494 329
rect 511 312 528 329
rect 545 312 562 329
rect 579 312 596 329
rect 613 312 630 329
rect 647 312 664 329
rect 681 312 767 329
rect 334 284 335 301
rect 352 284 353 301
rect 334 267 353 284
rect 551 285 573 293
rect 334 250 335 267
rect 352 251 353 267
rect 422 267 441 275
rect 422 262 423 267
rect 395 251 423 262
rect 352 250 423 251
rect 440 250 441 267
rect 334 240 441 250
rect 334 223 343 240
rect 360 233 441 240
rect 360 226 423 233
rect 360 223 364 226
rect 334 220 364 223
rect 334 215 360 220
rect 395 218 423 226
rect 334 198 335 215
rect 352 198 360 215
rect 422 216 423 218
rect 440 216 441 233
rect 422 207 441 216
rect 470 262 489 272
rect 470 245 471 262
rect 488 245 489 262
rect 470 228 489 245
rect 470 211 471 228
rect 488 211 489 228
rect 334 181 360 198
rect 470 185 489 211
rect 551 268 554 285
rect 571 268 573 285
rect 551 251 573 268
rect 551 234 554 251
rect 571 234 573 251
rect 551 206 573 234
rect 602 285 625 293
rect 602 268 607 285
rect 624 268 625 285
rect 602 254 625 268
rect 652 285 681 293
rect 669 268 681 285
rect 602 251 633 254
rect 602 234 607 251
rect 624 248 633 251
rect 602 231 616 234
rect 602 225 633 231
rect 652 251 681 268
rect 704 266 716 283
rect 733 266 745 283
rect 669 234 681 251
rect 710 239 740 266
rect 710 237 714 239
rect 735 237 740 239
rect 602 223 625 225
rect 551 189 635 206
rect 652 193 681 234
rect 704 220 714 237
rect 735 220 745 237
rect 710 218 714 220
rect 735 218 740 220
rect 710 193 740 218
rect 334 164 335 181
rect 352 164 360 181
rect 334 147 360 164
rect 439 182 489 185
rect 439 165 447 182
rect 464 165 489 182
rect 616 176 635 189
rect 439 162 489 165
rect 514 155 520 172
rect 537 155 571 172
rect 588 155 596 172
rect 616 167 638 176
rect 616 150 621 167
rect 616 147 638 150
rect 334 130 335 147
rect 352 130 360 147
rect 334 113 360 130
rect 334 96 335 113
rect 352 109 360 113
rect 396 136 442 144
rect 615 142 638 147
rect 396 119 423 136
rect 440 119 442 136
rect 396 117 442 119
rect 352 96 353 109
rect 334 86 353 96
rect 396 100 409 117
rect 426 100 442 117
rect 396 83 423 100
rect 440 83 442 100
rect 396 75 442 83
rect 469 130 490 142
rect 615 138 633 142
rect 469 113 471 130
rect 488 113 490 130
rect 469 96 490 113
rect 469 79 471 96
rect 488 79 490 96
rect 550 121 633 138
rect 550 109 572 121
rect 664 119 681 193
rect 704 176 716 193
rect 733 176 745 193
rect 550 92 554 109
rect 571 92 572 109
rect 651 104 681 119
rect 550 83 572 92
rect 603 95 625 103
rect 469 31 490 79
rect 603 78 607 95
rect 624 78 625 95
rect 603 70 625 78
rect 651 87 653 104
rect 670 87 681 104
rect 651 71 681 87
rect 0 14 80 31
rect 97 14 114 31
rect 131 14 148 31
rect 165 14 182 31
rect 199 14 216 31
rect 233 14 250 31
rect 267 14 284 31
rect 301 14 318 31
rect 335 14 352 31
rect 369 14 386 31
rect 403 14 420 31
rect 437 14 454 31
rect 471 14 488 31
rect 505 14 522 31
rect 539 14 556 31
rect 573 14 590 31
rect 607 14 624 31
rect 641 14 658 31
rect 675 14 767 31
<< viali >>
rect 80 605 97 622
rect 114 605 128 622
rect 128 605 131 622
rect 148 605 165 622
rect 182 605 199 622
rect 216 605 227 622
rect 227 605 233 622
rect 250 605 267 622
rect 284 605 292 622
rect 292 605 301 622
rect 318 605 335 622
rect 352 605 369 622
rect 386 605 391 622
rect 391 605 403 622
rect 420 605 437 622
rect 454 605 456 622
rect 456 605 471 622
rect 488 605 505 622
rect 522 605 539 622
rect 556 605 573 622
rect 590 605 607 622
rect 624 605 641 622
rect 658 605 675 622
rect 80 259 97 276
rect 98 206 115 223
rect 174 101 191 118
rect 287 130 304 141
rect 287 124 304 130
rect 494 312 511 329
rect 528 312 545 329
rect 562 312 579 329
rect 596 312 613 329
rect 630 312 647 329
rect 664 312 681 329
rect 343 223 360 240
rect 616 234 624 248
rect 624 234 633 248
rect 616 231 633 234
rect 714 237 735 239
rect 714 220 716 237
rect 716 220 733 237
rect 733 220 735 237
rect 714 218 735 220
rect 520 155 537 172
rect 409 100 426 117
rect 607 78 624 95
rect 80 14 97 31
rect 114 14 131 31
rect 148 14 165 31
rect 182 14 199 31
rect 216 14 233 31
rect 250 14 267 31
rect 284 14 301 31
rect 318 14 335 31
rect 352 14 369 31
rect 386 14 403 31
rect 420 14 437 31
rect 454 14 471 31
rect 488 14 505 31
rect 522 14 539 31
rect 556 14 573 31
rect 590 14 607 31
rect 624 14 641 31
rect 658 14 675 31
<< metal1 >>
rect 0 622 767 640
rect 0 605 80 622
rect 97 605 114 622
rect 131 605 148 622
rect 165 605 182 622
rect 199 605 216 622
rect 233 605 250 622
rect 267 605 284 622
rect 301 605 318 622
rect 335 605 352 622
rect 369 605 386 622
rect 403 605 420 622
rect 437 605 454 622
rect 471 605 488 622
rect 505 605 522 622
rect 539 605 556 622
rect 573 605 590 622
rect 607 605 624 622
rect 641 605 658 622
rect 675 605 767 622
rect 0 592 767 605
rect 0 329 767 344
rect 0 312 494 329
rect 511 312 528 329
rect 545 312 562 329
rect 579 312 596 329
rect 613 312 630 329
rect 647 312 664 329
rect 681 312 767 329
rect 0 296 767 312
rect 74 276 104 296
rect 74 259 80 276
rect 97 259 104 276
rect 74 253 104 259
rect 71 223 121 229
rect 71 206 98 223
rect 115 206 121 223
rect 71 201 121 206
rect 228 124 252 296
rect 334 246 369 249
rect 334 217 337 246
rect 366 217 369 246
rect 334 214 369 217
rect 513 176 545 179
rect 513 150 516 176
rect 542 150 545 176
rect 513 147 545 150
rect 168 118 252 124
rect 281 141 379 147
rect 281 124 287 141
rect 304 124 379 141
rect 281 123 379 124
rect 281 118 432 123
rect 168 101 174 118
rect 191 101 252 118
rect 168 95 252 101
rect 356 117 432 118
rect 356 100 409 117
rect 426 100 432 117
rect 356 94 432 100
rect 560 101 587 296
rect 610 248 741 254
rect 610 231 616 248
rect 633 239 741 248
rect 633 231 714 239
rect 610 225 714 231
rect 656 218 714 225
rect 735 218 741 239
rect 656 207 741 218
rect 560 95 627 101
rect 560 78 607 95
rect 624 78 627 95
rect 560 72 627 78
rect 656 48 686 207
rect 0 31 767 48
rect 0 14 80 31
rect 97 14 114 31
rect 131 14 148 31
rect 165 14 182 31
rect 199 14 216 31
rect 233 14 250 31
rect 267 14 284 31
rect 301 14 318 31
rect 335 14 352 31
rect 369 14 386 31
rect 403 14 420 31
rect 437 14 454 31
rect 471 14 488 31
rect 505 14 522 31
rect 539 14 556 31
rect 573 14 590 31
rect 607 14 624 31
rect 641 14 658 31
rect 675 14 767 31
rect 0 0 767 14
<< via1 >>
rect 337 240 366 246
rect 337 223 343 240
rect 343 223 360 240
rect 360 223 366 240
rect 337 217 366 223
rect 516 172 542 176
rect 516 155 520 172
rect 520 155 537 172
rect 537 155 542 172
rect 516 150 542 155
<< metal2 >>
rect 334 246 369 249
rect 334 217 337 246
rect 366 219 540 246
rect 366 217 369 219
rect 334 214 369 217
rect 514 179 540 219
rect 513 176 545 179
rect 513 150 516 176
rect 542 150 545 176
rect 513 147 545 150
<< labels >>
rlabel locali 664 149 681 166 1 Down
port 8 n signal output
rlabel locali 639 433 656 450 3 Up
port 7 n signal output
rlabel metal1 71 201 71 229 1 Clk2
port 9 n signal input
rlabel metal1 0 296 0 344 1 GND
port 11 n ground bidirectional
rlabel metal1 0 592 0 640 3 VDD
port 12 e power bidirectional
rlabel metal1 0 0 0 48 3 VDD
port 12 e power bidirectional
rlabel locali 87 146 114 173 1 Clk_Ref
port 3 n signal input
<< properties >>
string LEFclass CORE
string LEFsite unithddb1
<< end >>
