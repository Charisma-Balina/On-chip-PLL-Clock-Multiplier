* SKY130 Spice File.
*  Typical cell fet parameters
.param
+ sky130_fd_pr__special_nfet_latch__tox_mult = 1.000000    $ Units: meter
+ sky130_fd_pr__special_nfet_latch__lint_diff = 0.00    $ Units: meter
+ sky130_fd_pr__special_nfet_latch__wint_diff = 0.00    $ Units: meter
+ sky130_fd_pr__special_nfet_latch__deltal_diff = 0.00    $ Units: meter
+ sky130_fd_pr__special_nfet_latch__dlc_diff = 0.00    $ Units: meter
+ sky130_fd_pr__special_nfet_latch__dwc_diff = 0.00    $ Units: meter
+ sky130_fd_pr__special_nfet_latch__dvt0_diff = 0.00    $ Units: volt
+ sky130_fd_pr__special_nfet_latch__dvt1_diff = 0.00    $ Units: volt
+ sky130_fd_pr__special_nfet_latch__k3_diff = 0.0
+ sky130_fd_pr__special_nfet_latch__voff_diff_0 = 0.0
+ sky130_fd_pr__special_nfet_latch__kt1_diff_0 = 0.0
+ sky130_fd_pr__special_nfet_latch__rdsw_diff_0 = 0.0
+ sky130_fd_pr__special_nfet_latch__k2_diff_0 = 0.0
+ sky130_fd_pr__special_nfet_latch__u0_diff_0 = 0.000
+ sky130_fd_pr__special_nfet_latch__vth0_diff_0 = 0.0
+ sky130_fd_pr__special_nfet_latch__vsat_diff_0 = 0.0
+ sky130_fd_pr__special_nfet_latch__nfactor_diff_0 = 0.0
+ sky130_fd_pr__special_nfet_latch__ajunction_mult = 1.0
+ sky130_fd_pr__special_nfet_latch__pjunction_mult = 1.0
+ sky130_fd_pr__special_nfet_latch__overlap_mult = 1.0
+ sky130_fd_pr__special_nfet_latch__cit_diff = 0.00
+ sky130_fd_pr__special_nfet_latch__cdsc_diff = 0.00
+ sky130_fd_pr__special_nfet_latch__cdscb_diff = 0.00
+ sky130_fd_pr__special_nfet_latch__cdscd_diff = 0.00
+ sky130_fd_pr__special_nfet_latch__kt2_diff = 0.00
.param
+ sky130_fd_pr__special_nfet_pass__tox_mult = 1.000000    $ Units: meter
+ sky130_fd_pr__special_nfet_pass__lint_diff = 0.00    $ Units: meter
+ sky130_fd_pr__special_nfet_pass__wint_diff = 0.00    $ Units: meter
+ sky130_fd_pr__special_nfet_pass__deltal_diff = 0.00    $ Units: meter
+ sky130_fd_pr__special_nfet_pass__dlc_diff = 0.00    $ Units: meter
+ sky130_fd_pr__special_nfet_pass__dwc_diff = 0.00    $ Units: meter
+ sky130_fd_pr__special_nfet_pass__dvt0_diff = 0.00    $ Units: volt
+ sky130_fd_pr__special_nfet_pass__dvt1_diff = 0.00    $ Units: volt
+ sky130_fd_pr__special_nfet_pass__k3_diff = 0.0
+ sky130_fd_pr__special_nfet_pass__kt1_diff_0 = 0.0
+ sky130_fd_pr__special_nfet_pass__nfactor_diff_0 = 0.0
+ sky130_fd_pr__special_nfet_pass__vsat_diff_0 = 0.0
+ sky130_fd_pr__special_nfet_pass__k2_diff_0 = 0.0
+ sky130_fd_pr__special_nfet_pass__u0_diff_0 = -0.0
+ sky130_fd_pr__special_nfet_pass__vth0_diff_0 = 0.0
+ sky130_fd_pr__special_nfet_pass__rdsw_diff_0 = 0.0
+ sky130_fd_pr__special_nfet_pass__voff_diff_0 = 0.0
+ sky130_fd_pr__special_nfet_pass__ajunction_mult = 1.0
+ sky130_fd_pr__special_nfet_pass__pjunction_mult = 1.0
+ sky130_fd_pr__special_nfet_pass__overlap_mult = 1.0
+ sky130_fd_pr__special_nfet_pass__cit_diff = 0.00
+ sky130_fd_pr__special_nfet_pass__cdsc_diff = 0.00
+ sky130_fd_pr__special_nfet_pass__cdscb_diff = 0.00
+ sky130_fd_pr__special_nfet_pass__cdscd_diff = 0.00
+ sky130_fd_pr__special_nfet_pass__kt2_diff = 0.00
+ sky130_fd_pr__special_nfet_pass__kt1l_diff = 0.00
.param
+ sky130_fd_pr__special_pfet_pass__tox_mult = 1.0000    $ Units: meter
+ sky130_fd_pr__special_pfet_pass__lint_diff = 0.00    $ Units: meter
+ sky130_fd_pr__special_pfet_pass__wint_diff = 0.00    $ Units: meter
+ sky130_fd_pr__special_pfet_pass__dlc_diff = 0.00    $ Units: meter
+ sky130_fd_pr__special_pfet_pass__deltal_diff = 0.00    $ Units: meter
+ sky130_fd_pr__special_pfet_pass__deltaw_diff = 0.00    $ Units: meter
+ sky130_fd_pr__special_pfet_pass__dwc_diff = 0.00    $ Units: meter
+ sky130_fd_pr__special_pfet_pass__dvt0_diff = 0.00    $ Units: volt
+ sky130_fd_pr__special_pfet_pass__dvt1_diff = 0.00    $ Units: volt
+ sky130_fd_pr__special_pfet_pass__k3_diff = 0.0
+ sky130_fd_pr__special_pfet_pass__voff_diff_0 = 0.0
+ sky130_fd_pr__special_pfet_pass__kt1_diff_0 = 0.0
+ sky130_fd_pr__special_pfet_pass__vsat_diff_0 = 0.0
+ sky130_fd_pr__special_pfet_pass__vth0_diff_0 = 0.0
+ sky130_fd_pr__special_pfet_pass__nfactor_diff_0 = 0.0
+ sky130_fd_pr__special_pfet_pass__k2_diff_0 = 0.0
+ sky130_fd_pr__special_pfet_pass__u0_diff_0 = 0.0
+ sky130_fd_pr__special_pfet_pass__rdsw_diff_0 = 0.0
+ sky130_fd_pr__special_pfet_pass__ajunction_mult = 1.0
+ sky130_fd_pr__special_pfet_pass__pjunction_mult = 1.0
+ sky130_fd_pr__special_pfet_pass__overlap_mult = 1.00    $ Units: farad/meter
+ sky130_fd_pr__special_pfet_pass__cit_diff = 0.00
+ sky130_fd_pr__special_pfet_pass__cdsc_diff = 0.00
+ sky130_fd_pr__special_pfet_pass__cdscb_diff = 0.00
+ sky130_fd_pr__special_pfet_pass__cdscd_diff = 0.00
+ sky130_fd_pr__special_pfet_pass__kt2_diff = 0.00
+ sky130_fd_pr__special_pfet_pass__kt1l_diff = 0.00
* Typical Flash Nmos Pass Gate Parameters
.param
+ sky130_fd_pr__special_nfet_pass_flash__tox_mult = 1.00    $ Units: meter
+ sky130_fd_pr__special_nfet_pass_flash__lint_diff = 0.00    $ Units: meter
+ sky130_fd_pr__special_nfet_pass_flash__wint_diff = 0.00    $ Units: meter
+ sky130_fd_pr__special_nfet_pass_flash__dlc_diff = 0.00    $ Units: meter
+ sky130_fd_pr__special_nfet_pass_flash__dwc_diff = 0.00    $ Units: meter
+ sky130_fd_pr__special_nfet_pass_flash__dvt0_diff = 0.000   $ Units: volt
+ sky130_fd_pr__special_nfet_pass_flash__nlx_diff = 0.000   $ Units: volt
+ sky130_fd_pr__special_nfet_pass_flash__dvt1_diff = 0.00    $ Units: volt
+ sky130_fd_pr__special_nfet_pass_flash__dvt2_diff = 0.00    $ Units: volt
+ sky130_fd_pr__special_nfet_pass_flash__dvt0w_diff = 0.000   $ Units: volt
+ sky130_fd_pr__special_nfet_pass_flash__k3_diff = 000.0
+ sky130_fd_pr__special_nfet_pass_flash__k3b_diff = 000.0
+ sky130_fd_pr__special_nfet_pass_flash__ua_diff = 000.0
+ sky130_fd_pr__special_nfet_pass_flash__ub_diff = 000.0
+ sky130_fd_pr__special_nfet_pass_flash__uc_diff = 000.0
+ sky130_fd_pr__special_nfet_pass_flash__a0_diff = 000.0
+ sky130_fd_pr__special_nfet_pass_flash__ags_diff = 000.0
+ sky130_fd_pr__special_nfet_pass_flash__kt1_diff_0 = 0.0
+ sky130_fd_pr__special_nfet_pass_flash__nfactor_diff_0 = 0.0
+ sky130_fd_pr__special_nfet_pass_flash__voff_diff_0 = 0.0
+ sky130_fd_pr__special_nfet_pass_flash__k2_diff_0 = 0.0
+ sky130_fd_pr__special_nfet_pass_flash__u0_diff_0 = 0.0
+ sky130_fd_pr__special_nfet_pass_flash__vsat_diff_0 = 0.0
+ sky130_fd_pr__special_nfet_pass_flash__vth0_diff_0 = -0.0
+ sky130_fd_pr__special_nfet_pass_flash__kt1_diff_1 = 0.0
+ sky130_fd_pr__special_nfet_pass_flash__nfactor_diff_1 = 0.0
+ sky130_fd_pr__special_nfet_pass_flash__voff_diff_1 = 0.0
+ sky130_fd_pr__special_nfet_pass_flash__k2_diff_1 = 0.0
+ sky130_fd_pr__special_nfet_pass_flash__u0_diff_1 = 0.0
+ sky130_fd_pr__special_nfet_pass_flash__vsat_diff_1 = 0.0
+ sky130_fd_pr__special_nfet_pass_flash__vth0_diff_1 = -0.0
+ sky130_fd_pr__special_nfet_pass_flash__dwg_diff = 0.00    $ Units: volt
+ sky130_fd_pr__special_nfet_pass_flash__ajunction_mult = 1.0000    $ Units: farad/meter
+ sky130_fd_pr__special_nfet_pass_flash__pjunction_mult = 1.0000    $ Units: farad/meter
+ sky130_fd_pr__special_nfet_pass_flash__overlap_mult = 1.00      $ Units: farad/meter
+ sky130_fd_pr__special_nfet_pass_flash__cit_diff = 0.00
+ sky130_fd_pr__special_nfet_pass_flash__cdsc_diff = 0.00
+ sky130_fd_pr__special_nfet_pass_flash__cdscb_diff = 0.00
+ sky130_fd_pr__special_nfet_pass_flash__cdscd_diff = 0.00
+ sky130_fd_pr__special_nfet_pass_flash__kt2_diff = 0.00
+ sky130_fd_pr__special_nfet_pass_flash__kt1l_diff = 0.00
.include "../../../cells/special_nfet_latch/sky130_fd_pr__special_nfet_latch__mismatch.corner.spice"
.include "../../../cells/special_nfet_pass/sky130_fd_pr__special_nfet_pass__mismatch.corner.spice"
.include "../../../cells/special_nfet_pass_flash/sky130_fd_pr__special_nfet_pass_flash__mismatch.corner.spice"
.include "../../../cells/special_pfet_pass/sky130_fd_pr__special_pfet_pass__mismatch.corner.spice"
.include "../../../cells/special_nfet_pass_lvt/sky130_fd_pr__special_nfet_pass_lvt__wafer.corner.spice"
