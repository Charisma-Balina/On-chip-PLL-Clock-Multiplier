magic
tech sky130A
timestamp 1605998167
<< nwell >>
rect 12 467 2066 626
rect 12 436 816 467
rect 196 423 816 436
rect 230 408 816 423
rect 241 403 816 408
rect 1158 393 2066 467
rect 1158 389 1942 393
rect 1158 388 1288 389
rect 1158 358 1251 388
rect 60 117 315 168
rect 60 32 390 117
rect 1055 115 1139 160
rect 1055 31 1241 115
<< nmos >>
rect 860 360 902 375
rect 119 204 134 240
rect 243 204 258 240
rect 388 232 432 247
rect 462 232 942 247
rect 1054 233 1096 248
rect 462 176 1002 191
<< pmos >>
rect 248 565 2048 580
rect 172 516 216 531
rect 248 516 2048 531
rect 248 460 788 475
rect 1185 409 1227 424
rect 119 73 134 145
rect 243 74 258 146
rect 1073 94 1115 109
<< ndiff >>
rect 860 400 902 408
rect 860 383 873 400
rect 890 383 902 400
rect 860 375 902 383
rect 860 352 902 360
rect 860 335 873 352
rect 890 335 902 352
rect 860 327 902 335
rect 388 272 432 280
rect 388 255 401 272
rect 418 255 432 272
rect 388 247 432 255
rect 462 272 942 280
rect 462 255 466 272
rect 483 255 500 272
rect 517 255 534 272
rect 551 255 568 272
rect 585 255 602 272
rect 619 255 636 272
rect 653 255 670 272
rect 687 255 704 272
rect 721 255 738 272
rect 755 255 772 272
rect 789 255 806 272
rect 823 255 840 272
rect 857 255 874 272
rect 891 255 908 272
rect 925 255 942 272
rect 462 247 942 255
rect 1054 273 1096 281
rect 1054 256 1070 273
rect 1087 256 1096 273
rect 1054 248 1096 256
rect 87 230 119 240
rect 87 213 94 230
rect 111 213 119 230
rect 87 204 119 213
rect 134 230 167 240
rect 134 213 142 230
rect 159 213 167 230
rect 134 204 167 213
rect 211 230 243 240
rect 211 213 218 230
rect 235 213 243 230
rect 211 204 243 213
rect 258 230 291 240
rect 258 213 266 230
rect 283 213 291 230
rect 258 204 291 213
rect 388 224 432 232
rect 388 207 401 224
rect 418 207 432 224
rect 388 199 432 207
rect 462 224 942 232
rect 462 216 1002 224
rect 462 199 470 216
rect 487 199 504 216
rect 521 199 538 216
rect 555 199 572 216
rect 589 199 606 216
rect 623 199 640 216
rect 657 199 674 216
rect 691 199 708 216
rect 725 199 742 216
rect 759 199 776 216
rect 793 199 810 216
rect 827 199 844 216
rect 861 199 878 216
rect 895 199 912 216
rect 929 199 946 216
rect 963 199 1002 216
rect 1054 221 1096 233
rect 1054 204 1067 221
rect 1084 204 1096 221
rect 1054 200 1096 204
rect 462 191 1002 199
rect 462 168 1002 176
rect 462 151 470 168
rect 487 151 504 168
rect 521 151 538 168
rect 555 151 572 168
rect 589 151 606 168
rect 623 151 640 168
rect 657 151 674 168
rect 691 151 708 168
rect 725 151 742 168
rect 759 151 776 168
rect 793 151 810 168
rect 827 151 844 168
rect 861 151 878 168
rect 895 151 912 168
rect 929 151 946 168
rect 963 151 1002 168
rect 462 143 1002 151
<< pdiff >>
rect 248 603 2048 608
rect 248 586 257 603
rect 274 586 291 603
rect 308 586 325 603
rect 342 586 359 603
rect 376 586 393 603
rect 410 586 427 603
rect 444 586 461 603
rect 478 586 495 603
rect 512 586 529 603
rect 546 586 563 603
rect 580 586 597 603
rect 614 586 631 603
rect 648 586 665 603
rect 682 586 699 603
rect 716 586 733 603
rect 750 586 767 603
rect 784 586 801 603
rect 818 586 835 603
rect 852 586 869 603
rect 886 586 903 603
rect 920 586 937 603
rect 954 586 971 603
rect 988 586 1005 603
rect 1022 586 1039 603
rect 1056 586 1073 603
rect 1090 586 1107 603
rect 1124 586 1141 603
rect 1158 586 1175 603
rect 1192 586 1209 603
rect 1226 586 1243 603
rect 1260 586 1277 603
rect 1294 586 1311 603
rect 1328 586 1345 603
rect 1362 586 1379 603
rect 1396 586 1413 603
rect 1430 586 1447 603
rect 1464 586 1481 603
rect 1498 586 1515 603
rect 1532 586 1549 603
rect 1566 586 1583 603
rect 1600 586 1617 603
rect 1634 586 1651 603
rect 1668 586 1685 603
rect 1702 586 1719 603
rect 1736 586 1753 603
rect 1770 586 1787 603
rect 1804 586 1821 603
rect 1838 586 1855 603
rect 1872 586 1889 603
rect 1906 586 1923 603
rect 1940 586 1957 603
rect 1974 586 1991 603
rect 2008 586 2048 603
rect 248 580 2048 586
rect 172 557 216 565
rect 172 540 185 557
rect 202 540 216 557
rect 172 531 216 540
rect 248 557 2048 565
rect 248 540 257 557
rect 274 540 291 557
rect 308 540 325 557
rect 342 540 359 557
rect 376 540 393 557
rect 410 540 427 557
rect 444 540 461 557
rect 478 540 495 557
rect 512 540 529 557
rect 546 540 563 557
rect 580 540 597 557
rect 614 540 631 557
rect 648 540 665 557
rect 682 540 699 557
rect 716 540 733 557
rect 750 540 767 557
rect 784 540 801 557
rect 818 540 835 557
rect 852 540 869 557
rect 886 540 903 557
rect 920 540 937 557
rect 954 540 971 557
rect 988 540 1005 557
rect 1022 540 1039 557
rect 1056 540 1073 557
rect 1090 540 1107 557
rect 1124 540 1141 557
rect 1158 540 1175 557
rect 1192 540 1209 557
rect 1226 540 1243 557
rect 1260 540 1277 557
rect 1294 540 1311 557
rect 1328 540 1345 557
rect 1362 540 1379 557
rect 1396 540 1413 557
rect 1430 540 1447 557
rect 1464 540 1481 557
rect 1498 540 1515 557
rect 1532 540 1549 557
rect 1566 540 1583 557
rect 1600 540 1617 557
rect 1634 540 1651 557
rect 1668 540 1685 557
rect 1702 540 1719 557
rect 1736 540 1753 557
rect 1770 540 1787 557
rect 1804 540 1821 557
rect 1838 540 1855 557
rect 1872 540 1889 557
rect 1906 540 1923 557
rect 1940 540 1957 557
rect 1974 540 1991 557
rect 2008 540 2048 557
rect 248 531 2048 540
rect 172 508 216 516
rect 172 491 186 508
rect 203 491 216 508
rect 172 483 216 491
rect 248 508 2048 516
rect 248 491 257 508
rect 274 491 291 508
rect 308 491 325 508
rect 342 491 359 508
rect 376 491 393 508
rect 410 491 427 508
rect 444 491 461 508
rect 478 491 495 508
rect 512 491 529 508
rect 546 491 563 508
rect 580 491 597 508
rect 614 491 631 508
rect 648 491 665 508
rect 682 491 699 508
rect 716 491 733 508
rect 750 491 767 508
rect 784 491 801 508
rect 818 491 835 508
rect 852 491 869 508
rect 886 491 903 508
rect 920 491 937 508
rect 954 491 971 508
rect 988 491 1005 508
rect 1022 491 1039 508
rect 1056 491 1073 508
rect 1090 491 1107 508
rect 1124 491 1141 508
rect 1158 491 1175 508
rect 1192 491 1209 508
rect 1226 491 1243 508
rect 1260 491 1277 508
rect 1294 491 1311 508
rect 1328 491 1345 508
rect 1362 491 1379 508
rect 1396 491 1413 508
rect 1430 491 1447 508
rect 1464 491 1481 508
rect 1498 491 1515 508
rect 1532 491 1549 508
rect 1566 491 1583 508
rect 1600 491 1617 508
rect 1634 491 1651 508
rect 1668 491 1685 508
rect 1702 491 1719 508
rect 1736 491 1753 508
rect 1770 491 1787 508
rect 1804 491 1821 508
rect 1838 491 1855 508
rect 1872 491 1889 508
rect 1906 491 1923 508
rect 1940 491 1957 508
rect 1974 491 1991 508
rect 2008 491 2048 508
rect 248 485 2048 491
rect 248 475 788 485
rect 248 452 788 460
rect 248 435 257 452
rect 274 435 291 452
rect 308 435 325 452
rect 342 435 359 452
rect 376 435 393 452
rect 410 435 427 452
rect 444 435 461 452
rect 478 435 495 452
rect 512 435 529 452
rect 546 435 563 452
rect 580 435 597 452
rect 614 435 631 452
rect 648 435 665 452
rect 682 435 699 452
rect 716 435 733 452
rect 750 435 788 452
rect 248 427 788 435
rect 1185 449 1227 457
rect 1185 432 1198 449
rect 1215 432 1227 449
rect 1185 424 1227 432
rect 1185 401 1227 409
rect 1185 384 1194 401
rect 1211 384 1227 401
rect 1185 376 1227 384
rect 86 128 119 145
rect 86 111 94 128
rect 111 111 119 128
rect 86 94 119 111
rect 86 77 94 94
rect 111 77 119 94
rect 86 73 119 77
rect 134 141 167 145
rect 134 124 142 141
rect 159 124 167 141
rect 134 107 167 124
rect 134 90 142 107
rect 159 90 167 107
rect 134 73 167 90
rect 210 129 243 146
rect 210 112 218 129
rect 235 112 243 129
rect 210 95 243 112
rect 210 78 218 95
rect 235 78 243 95
rect 210 74 243 78
rect 258 142 291 146
rect 258 125 266 142
rect 283 125 291 142
rect 258 108 291 125
rect 1073 134 1115 142
rect 258 91 266 108
rect 283 91 291 108
rect 258 74 291 91
rect 1073 117 1086 134
rect 1103 117 1115 134
rect 1073 109 1115 117
rect 1073 86 1115 94
rect 1073 69 1086 86
rect 1103 69 1115 86
rect 1073 61 1115 69
<< ndiffc >>
rect 873 383 890 400
rect 873 335 890 352
rect 401 255 418 272
rect 466 255 483 272
rect 500 255 517 272
rect 534 255 551 272
rect 568 255 585 272
rect 602 255 619 272
rect 636 255 653 272
rect 670 255 687 272
rect 704 255 721 272
rect 738 255 755 272
rect 772 255 789 272
rect 806 255 823 272
rect 840 255 857 272
rect 874 255 891 272
rect 908 255 925 272
rect 1070 256 1087 273
rect 94 213 111 230
rect 142 213 159 230
rect 218 213 235 230
rect 266 213 283 230
rect 401 207 418 224
rect 470 199 487 216
rect 504 199 521 216
rect 538 199 555 216
rect 572 199 589 216
rect 606 199 623 216
rect 640 199 657 216
rect 674 199 691 216
rect 708 199 725 216
rect 742 199 759 216
rect 776 199 793 216
rect 810 199 827 216
rect 844 199 861 216
rect 878 199 895 216
rect 912 199 929 216
rect 946 199 963 216
rect 1067 204 1084 221
rect 470 151 487 168
rect 504 151 521 168
rect 538 151 555 168
rect 572 151 589 168
rect 606 151 623 168
rect 640 151 657 168
rect 674 151 691 168
rect 708 151 725 168
rect 742 151 759 168
rect 776 151 793 168
rect 810 151 827 168
rect 844 151 861 168
rect 878 151 895 168
rect 912 151 929 168
rect 946 151 963 168
<< pdiffc >>
rect 257 586 274 603
rect 291 586 308 603
rect 325 586 342 603
rect 359 586 376 603
rect 393 586 410 603
rect 427 586 444 603
rect 461 586 478 603
rect 495 586 512 603
rect 529 586 546 603
rect 563 586 580 603
rect 597 586 614 603
rect 631 586 648 603
rect 665 586 682 603
rect 699 586 716 603
rect 733 586 750 603
rect 767 586 784 603
rect 801 586 818 603
rect 835 586 852 603
rect 869 586 886 603
rect 903 586 920 603
rect 937 586 954 603
rect 971 586 988 603
rect 1005 586 1022 603
rect 1039 586 1056 603
rect 1073 586 1090 603
rect 1107 586 1124 603
rect 1141 586 1158 603
rect 1175 586 1192 603
rect 1209 586 1226 603
rect 1243 586 1260 603
rect 1277 586 1294 603
rect 1311 586 1328 603
rect 1345 586 1362 603
rect 1379 586 1396 603
rect 1413 586 1430 603
rect 1447 586 1464 603
rect 1481 586 1498 603
rect 1515 586 1532 603
rect 1549 586 1566 603
rect 1583 586 1600 603
rect 1617 586 1634 603
rect 1651 586 1668 603
rect 1685 586 1702 603
rect 1719 586 1736 603
rect 1753 586 1770 603
rect 1787 586 1804 603
rect 1821 586 1838 603
rect 1855 586 1872 603
rect 1889 586 1906 603
rect 1923 586 1940 603
rect 1957 586 1974 603
rect 1991 586 2008 603
rect 185 540 202 557
rect 257 540 274 557
rect 291 540 308 557
rect 325 540 342 557
rect 359 540 376 557
rect 393 540 410 557
rect 427 540 444 557
rect 461 540 478 557
rect 495 540 512 557
rect 529 540 546 557
rect 563 540 580 557
rect 597 540 614 557
rect 631 540 648 557
rect 665 540 682 557
rect 699 540 716 557
rect 733 540 750 557
rect 767 540 784 557
rect 801 540 818 557
rect 835 540 852 557
rect 869 540 886 557
rect 903 540 920 557
rect 937 540 954 557
rect 971 540 988 557
rect 1005 540 1022 557
rect 1039 540 1056 557
rect 1073 540 1090 557
rect 1107 540 1124 557
rect 1141 540 1158 557
rect 1175 540 1192 557
rect 1209 540 1226 557
rect 1243 540 1260 557
rect 1277 540 1294 557
rect 1311 540 1328 557
rect 1345 540 1362 557
rect 1379 540 1396 557
rect 1413 540 1430 557
rect 1447 540 1464 557
rect 1481 540 1498 557
rect 1515 540 1532 557
rect 1549 540 1566 557
rect 1583 540 1600 557
rect 1617 540 1634 557
rect 1651 540 1668 557
rect 1685 540 1702 557
rect 1719 540 1736 557
rect 1753 540 1770 557
rect 1787 540 1804 557
rect 1821 540 1838 557
rect 1855 540 1872 557
rect 1889 540 1906 557
rect 1923 540 1940 557
rect 1957 540 1974 557
rect 1991 540 2008 557
rect 186 491 203 508
rect 257 491 274 508
rect 291 491 308 508
rect 325 491 342 508
rect 359 491 376 508
rect 393 491 410 508
rect 427 491 444 508
rect 461 491 478 508
rect 495 491 512 508
rect 529 491 546 508
rect 563 491 580 508
rect 597 491 614 508
rect 631 491 648 508
rect 665 491 682 508
rect 699 491 716 508
rect 733 491 750 508
rect 767 491 784 508
rect 801 491 818 508
rect 835 491 852 508
rect 869 491 886 508
rect 903 491 920 508
rect 937 491 954 508
rect 971 491 988 508
rect 1005 491 1022 508
rect 1039 491 1056 508
rect 1073 491 1090 508
rect 1107 491 1124 508
rect 1141 491 1158 508
rect 1175 491 1192 508
rect 1209 491 1226 508
rect 1243 491 1260 508
rect 1277 491 1294 508
rect 1311 491 1328 508
rect 1345 491 1362 508
rect 1379 491 1396 508
rect 1413 491 1430 508
rect 1447 491 1464 508
rect 1481 491 1498 508
rect 1515 491 1532 508
rect 1549 491 1566 508
rect 1583 491 1600 508
rect 1617 491 1634 508
rect 1651 491 1668 508
rect 1685 491 1702 508
rect 1719 491 1736 508
rect 1753 491 1770 508
rect 1787 491 1804 508
rect 1821 491 1838 508
rect 1855 491 1872 508
rect 1889 491 1906 508
rect 1923 491 1940 508
rect 1957 491 1974 508
rect 1991 491 2008 508
rect 257 435 274 452
rect 291 435 308 452
rect 325 435 342 452
rect 359 435 376 452
rect 393 435 410 452
rect 427 435 444 452
rect 461 435 478 452
rect 495 435 512 452
rect 529 435 546 452
rect 563 435 580 452
rect 597 435 614 452
rect 631 435 648 452
rect 665 435 682 452
rect 699 435 716 452
rect 733 435 750 452
rect 1198 432 1215 449
rect 1194 384 1211 401
rect 94 111 111 128
rect 94 77 111 94
rect 142 124 159 141
rect 142 90 159 107
rect 218 112 235 129
rect 218 78 235 95
rect 266 125 283 142
rect 266 91 283 108
rect 1086 117 1103 134
rect 1086 69 1103 86
<< psubdiff >>
rect 145 332 157 349
rect 174 332 186 349
rect 227 332 239 349
rect 256 332 268 349
rect 309 332 321 349
rect 338 332 350 349
rect 391 332 403 349
rect 420 332 432 349
rect 473 332 485 349
rect 502 332 514 349
rect 555 332 567 349
rect 584 332 596 349
rect 1223 287 1235 304
rect 1252 287 1264 304
rect 1305 287 1317 304
rect 1334 287 1346 304
rect 1387 287 1399 304
rect 1416 287 1428 304
rect 1469 287 1481 304
rect 1498 287 1510 304
rect 1551 287 1563 304
rect 1580 287 1592 304
rect 1633 287 1645 304
rect 1662 287 1674 304
rect 1711 287 1723 304
rect 1740 287 1752 304
rect 1793 287 1805 304
rect 1822 287 1834 304
rect 1875 287 1887 304
rect 1904 287 1916 304
<< nsubdiff >>
rect 1339 422 1351 439
rect 1368 422 1380 439
rect 1421 422 1433 439
rect 1450 422 1462 439
rect 1503 422 1515 439
rect 1532 422 1544 439
rect 1585 422 1597 439
rect 1614 422 1626 439
rect 1667 422 1679 439
rect 1696 422 1708 439
rect 1749 422 1761 439
rect 1778 422 1790 439
rect 1831 422 1843 439
rect 1860 422 1872 439
rect 1913 422 1925 439
rect 1942 422 1954 439
rect 331 50 343 67
rect 360 50 372 67
rect 1168 61 1180 78
rect 1197 61 1209 78
<< psubdiffcont >>
rect 157 332 174 349
rect 239 332 256 349
rect 321 332 338 349
rect 403 332 420 349
rect 485 332 502 349
rect 567 332 584 349
rect 1235 287 1252 304
rect 1317 287 1334 304
rect 1399 287 1416 304
rect 1481 287 1498 304
rect 1563 287 1580 304
rect 1645 287 1662 304
rect 1723 287 1740 304
rect 1805 287 1822 304
rect 1887 287 1904 304
<< nsubdiffcont >>
rect 1351 422 1368 439
rect 1433 422 1450 439
rect 1515 422 1532 439
rect 1597 422 1614 439
rect 1679 422 1696 439
rect 1761 422 1778 439
rect 1843 422 1860 439
rect 1925 422 1942 439
rect 343 50 360 67
rect 1180 61 1197 78
<< poly >>
rect 54 580 240 598
rect 54 509 73 580
rect 225 565 248 580
rect 2048 565 2061 580
rect 137 516 172 531
rect 216 516 248 531
rect 2048 516 2061 531
rect 130 513 152 516
rect 54 501 98 509
rect 54 484 69 501
rect 86 484 98 501
rect 125 508 152 513
rect 125 491 130 508
rect 147 491 152 508
rect 125 486 152 491
rect 54 477 98 484
rect 130 483 152 486
rect 219 460 248 475
rect 788 460 801 475
rect 219 433 236 460
rect 196 428 236 433
rect 196 411 204 428
rect 221 411 236 428
rect 196 406 236 411
rect 1122 425 1171 430
rect 1122 408 1130 425
rect 1147 424 1171 425
rect 1147 409 1185 424
rect 1227 409 1240 424
rect 1147 408 1171 409
rect 1122 403 1171 408
rect 798 376 825 384
rect 798 359 803 376
rect 820 375 825 376
rect 820 360 860 375
rect 902 360 915 375
rect 820 359 825 360
rect 798 351 825 359
rect 119 240 134 253
rect 243 240 258 253
rect 1002 274 1035 280
rect 1002 257 1010 274
rect 1027 257 1035 274
rect 1002 252 1035 257
rect 1017 248 1035 252
rect 352 232 388 247
rect 432 232 462 247
rect 942 232 957 247
rect 1017 233 1054 248
rect 1096 233 1109 248
rect 345 229 367 232
rect 340 224 367 229
rect 340 207 345 224
rect 362 207 367 224
rect 119 188 134 204
rect 243 188 258 204
rect 340 202 367 207
rect 345 199 367 202
rect 70 183 134 188
rect 70 166 78 183
rect 95 166 134 183
rect 70 161 134 166
rect 194 183 258 188
rect 194 166 202 183
rect 219 166 258 183
rect 425 176 462 191
rect 1002 176 1015 191
rect 425 171 449 176
rect 194 161 258 166
rect 119 145 134 161
rect 243 146 258 161
rect 400 166 449 171
rect 400 146 408 166
rect 429 146 449 166
rect 400 141 449 146
rect 1016 110 1043 118
rect 1016 93 1021 110
rect 1038 109 1043 110
rect 1038 94 1073 109
rect 1115 94 1128 109
rect 1038 93 1043 94
rect 1016 85 1043 93
rect 119 60 134 73
rect 243 61 258 74
<< polycont >>
rect 69 484 86 501
rect 130 491 147 508
rect 204 411 221 428
rect 1130 408 1147 425
rect 803 359 820 376
rect 1010 257 1027 274
rect 345 207 362 224
rect 78 166 95 183
rect 202 166 219 183
rect 408 146 429 166
rect 1021 93 1038 110
<< locali >>
rect 0 607 21 624
rect 38 607 55 624
rect 72 607 89 624
rect 106 607 123 624
rect 140 607 157 624
rect 174 607 191 624
rect 208 607 225 624
rect 242 607 259 624
rect 276 607 293 624
rect 310 607 327 624
rect 344 607 361 624
rect 378 607 395 624
rect 412 607 429 624
rect 446 607 463 624
rect 480 607 497 624
rect 514 607 531 624
rect 548 607 565 624
rect 582 607 599 624
rect 616 607 633 624
rect 650 607 667 624
rect 684 607 701 624
rect 718 607 735 624
rect 752 607 769 624
rect 786 607 803 624
rect 820 607 837 624
rect 854 607 871 624
rect 888 607 905 624
rect 922 607 939 624
rect 956 607 973 624
rect 990 607 1007 624
rect 1024 607 1041 624
rect 1058 607 1075 624
rect 1092 607 1109 624
rect 1126 607 1143 624
rect 1160 607 1177 624
rect 1194 607 1211 624
rect 1228 607 1245 624
rect 1262 607 1279 624
rect 1296 607 1313 624
rect 1330 607 1347 624
rect 1364 607 1381 624
rect 1398 607 1415 624
rect 1432 607 1449 624
rect 1466 607 1483 624
rect 1500 607 1517 624
rect 1534 607 1551 624
rect 1568 607 1585 624
rect 1602 607 1619 624
rect 1636 607 1653 624
rect 1670 607 1687 624
rect 1704 607 1721 624
rect 1738 607 1755 624
rect 1772 607 1789 624
rect 1806 607 1823 624
rect 1840 607 1857 624
rect 1874 607 1891 624
rect 1908 607 1925 624
rect 1942 607 1959 624
rect 1976 607 1993 624
rect 2010 607 2027 624
rect 2044 607 2066 624
rect 248 603 2048 607
rect 248 586 257 603
rect 274 586 291 603
rect 308 586 325 603
rect 342 586 359 603
rect 376 586 393 603
rect 410 586 427 603
rect 444 586 461 603
rect 478 586 495 603
rect 512 586 529 603
rect 546 586 563 603
rect 580 586 597 603
rect 614 586 631 603
rect 648 586 665 603
rect 682 586 699 603
rect 716 586 733 603
rect 750 586 767 603
rect 784 586 801 603
rect 818 586 835 603
rect 852 586 869 603
rect 886 586 903 603
rect 920 586 937 603
rect 954 586 971 603
rect 988 586 1005 603
rect 1022 586 1039 603
rect 1056 586 1073 603
rect 1090 586 1107 603
rect 1124 586 1141 603
rect 1158 586 1175 603
rect 1192 586 1209 603
rect 1226 586 1243 603
rect 1260 586 1277 603
rect 1294 586 1311 603
rect 1328 586 1345 603
rect 1362 586 1379 603
rect 1396 586 1413 603
rect 1430 586 1447 603
rect 1464 586 1481 603
rect 1498 586 1515 603
rect 1532 586 1549 603
rect 1566 586 1583 603
rect 1600 586 1617 603
rect 1634 586 1651 603
rect 1668 586 1685 603
rect 1702 586 1719 603
rect 1736 586 1753 603
rect 1770 586 1787 603
rect 1804 586 1821 603
rect 1838 586 1855 603
rect 1872 586 1889 603
rect 1906 586 1923 603
rect 1940 586 1957 603
rect 1974 586 1991 603
rect 2008 586 2048 603
rect 248 585 2048 586
rect 172 557 2048 558
rect 172 540 185 557
rect 202 540 257 557
rect 274 540 291 557
rect 308 540 325 557
rect 342 540 359 557
rect 376 540 393 557
rect 410 540 427 557
rect 444 540 461 557
rect 478 540 495 557
rect 512 540 529 557
rect 546 540 563 557
rect 580 540 597 557
rect 614 540 631 557
rect 648 540 665 557
rect 682 540 699 557
rect 716 540 733 557
rect 750 540 767 557
rect 784 540 801 557
rect 818 540 835 557
rect 852 540 869 557
rect 886 540 903 557
rect 920 540 937 557
rect 954 540 971 557
rect 988 540 1005 557
rect 1022 540 1039 557
rect 1056 540 1073 557
rect 1090 540 1107 557
rect 1124 540 1141 557
rect 1158 540 1175 557
rect 1192 540 1209 557
rect 1226 540 1243 557
rect 1260 540 1277 557
rect 1298 540 1311 557
rect 1332 540 1345 557
rect 1362 540 1379 557
rect 1396 540 1413 557
rect 1430 540 1447 557
rect 1464 540 1481 557
rect 1498 540 1515 557
rect 1532 540 1549 557
rect 1566 540 1583 557
rect 1600 540 1617 557
rect 1634 540 1651 557
rect 1668 540 1685 557
rect 1702 540 1719 557
rect 1736 540 1753 557
rect 1770 540 1787 557
rect 1804 540 1821 557
rect 1838 540 1855 557
rect 1872 540 1889 557
rect 1906 540 1923 557
rect 1940 540 1957 557
rect 1974 540 1991 557
rect 2008 540 2048 557
rect 172 539 2048 540
rect 837 534 875 539
rect 963 534 1001 539
rect 1187 534 1225 539
rect 122 508 216 509
rect 51 501 96 505
rect 51 484 69 501
rect 86 484 96 501
rect 122 491 130 508
rect 147 491 186 508
rect 203 491 216 508
rect 122 490 216 491
rect 248 508 2048 509
rect 248 491 257 508
rect 274 491 291 508
rect 308 491 325 508
rect 342 491 359 508
rect 376 491 393 508
rect 410 491 427 508
rect 444 491 461 508
rect 478 491 495 508
rect 512 491 529 508
rect 546 491 563 508
rect 580 491 597 508
rect 614 491 631 508
rect 648 491 665 508
rect 682 491 699 508
rect 716 491 733 508
rect 750 491 767 508
rect 784 491 801 508
rect 818 491 835 508
rect 852 491 869 508
rect 886 491 903 508
rect 920 491 937 508
rect 954 491 971 508
rect 988 491 1005 508
rect 1022 491 1039 508
rect 1056 491 1073 508
rect 1090 491 1107 508
rect 1124 491 1141 508
rect 1158 491 1175 508
rect 1192 491 1209 508
rect 1226 491 1243 508
rect 1260 491 1277 508
rect 1294 491 1311 508
rect 1328 491 1345 508
rect 1362 491 1379 508
rect 1396 491 1413 508
rect 1430 491 1447 508
rect 1464 491 1481 508
rect 1498 491 1515 508
rect 1532 491 1549 508
rect 1566 491 1583 508
rect 1600 491 1617 508
rect 1634 491 1651 508
rect 1668 491 1685 508
rect 1702 491 1719 508
rect 1736 491 1753 508
rect 1770 491 1787 508
rect 1804 491 1821 508
rect 1838 491 1855 508
rect 1872 491 1889 508
rect 1906 491 1923 508
rect 1940 491 1957 508
rect 1974 491 1991 508
rect 2008 491 2048 508
rect 248 490 2048 491
rect 837 485 875 490
rect 963 485 1001 490
rect 51 481 96 484
rect 204 428 221 436
rect 248 435 257 452
rect 274 435 291 452
rect 308 435 325 452
rect 342 435 359 452
rect 376 435 393 452
rect 410 435 427 452
rect 444 435 461 452
rect 478 435 495 452
rect 512 435 529 452
rect 546 435 563 452
rect 580 435 597 452
rect 614 435 631 452
rect 648 435 665 452
rect 682 435 699 452
rect 716 435 733 452
rect 750 435 902 452
rect 1187 450 1225 490
rect 204 403 221 411
rect 799 376 824 435
rect 843 430 902 435
rect 1185 449 1227 450
rect 1185 432 1198 449
rect 1215 432 1227 449
rect 1185 431 1227 432
rect 1338 439 2015 441
rect 848 425 902 430
rect 855 419 902 425
rect 860 400 902 419
rect 1122 408 1130 425
rect 1147 408 1155 425
rect 1338 422 1351 439
rect 1368 422 1433 439
rect 1450 422 1515 439
rect 1532 422 1597 439
rect 1614 422 1679 439
rect 1696 422 1761 439
rect 1778 422 1843 439
rect 1860 422 1882 439
rect 1899 422 1925 439
rect 1942 422 2015 439
rect 1338 420 2015 422
rect 860 383 873 400
rect 890 383 902 400
rect 1185 401 2066 402
rect 1185 387 1194 401
rect 1061 384 1194 387
rect 1211 384 2066 401
rect 795 359 803 376
rect 820 359 828 376
rect 130 349 637 355
rect 130 332 157 349
rect 174 332 239 349
rect 256 332 321 349
rect 338 332 403 349
rect 420 332 485 349
rect 502 332 567 349
rect 584 332 637 349
rect 130 327 637 332
rect 860 335 873 352
rect 890 335 902 352
rect 860 327 902 335
rect 1061 349 2066 384
rect 1061 348 1196 349
rect 1 310 21 327
rect 38 310 55 327
rect 72 310 89 327
rect 106 310 123 327
rect 140 310 157 327
rect 174 310 191 327
rect 208 310 225 327
rect 242 310 259 327
rect 276 310 293 327
rect 310 310 327 327
rect 344 310 361 327
rect 378 310 395 327
rect 412 310 429 327
rect 446 310 463 327
rect 480 310 497 327
rect 514 310 531 327
rect 548 310 565 327
rect 582 310 599 327
rect 616 310 633 327
rect 650 310 667 327
rect 684 310 701 327
rect 718 310 735 327
rect 752 310 769 327
rect 786 310 803 327
rect 820 310 837 327
rect 854 310 871 327
rect 888 310 905 327
rect 922 310 939 327
rect 956 310 973 327
rect 990 310 1007 327
rect 1024 310 1041 327
rect 93 230 112 310
rect 93 213 94 230
rect 111 213 112 230
rect 93 204 112 213
rect 141 271 167 276
rect 141 254 146 271
rect 163 254 167 271
rect 141 250 167 254
rect 141 230 160 250
rect 141 213 142 230
rect 159 213 160 230
rect 70 166 78 183
rect 95 166 103 183
rect 93 128 112 145
rect 93 111 94 128
rect 111 111 112 128
rect 93 94 112 111
rect 93 77 94 94
rect 111 77 112 94
rect 93 69 112 77
rect 141 141 160 213
rect 217 230 236 310
rect 401 273 925 310
rect 1010 274 1027 282
rect 401 272 942 273
rect 388 255 401 272
rect 418 255 466 272
rect 483 255 500 272
rect 517 255 534 272
rect 551 255 568 272
rect 585 255 602 272
rect 619 255 636 272
rect 653 255 670 272
rect 687 255 704 272
rect 721 255 738 272
rect 755 255 772 272
rect 789 255 806 272
rect 823 255 840 272
rect 857 255 874 272
rect 891 255 908 272
rect 925 255 942 272
rect 462 254 942 255
rect 1061 273 1096 348
rect 1114 310 1143 327
rect 1160 310 1177 327
rect 1194 310 1211 327
rect 1228 310 1245 327
rect 1262 310 1279 327
rect 1296 310 1313 327
rect 1330 310 1347 327
rect 1364 310 1381 327
rect 1398 310 1415 327
rect 1432 310 1449 327
rect 1466 310 1483 327
rect 1500 310 1517 327
rect 1534 310 1551 327
rect 1568 310 1585 327
rect 1602 310 1619 327
rect 1636 310 1653 327
rect 1670 310 1687 327
rect 1704 310 1721 327
rect 1738 310 1755 327
rect 1772 310 1789 327
rect 1806 310 1823 327
rect 1840 310 1857 327
rect 1874 310 1891 327
rect 1908 310 1925 327
rect 1942 310 1959 327
rect 1976 310 1993 327
rect 2010 310 2066 327
rect 1208 304 1957 310
rect 1208 287 1235 304
rect 1252 287 1317 304
rect 1334 287 1399 304
rect 1416 287 1481 304
rect 1498 287 1563 304
rect 1580 287 1645 304
rect 1662 287 1723 304
rect 1740 287 1805 304
rect 1822 287 1887 304
rect 1904 287 1957 304
rect 1208 282 1957 287
rect 1010 249 1027 257
rect 1054 256 1070 273
rect 1087 256 1096 273
rect 217 213 218 230
rect 235 213 236 230
rect 217 204 236 213
rect 265 230 284 240
rect 265 213 266 230
rect 283 213 284 230
rect 194 166 202 183
rect 219 166 227 183
rect 265 174 284 213
rect 337 224 432 225
rect 337 207 345 224
rect 362 207 401 224
rect 418 207 432 224
rect 1054 222 1096 225
rect 999 221 1096 222
rect 999 217 1067 221
rect 337 206 432 207
rect 462 216 1067 217
rect 462 199 470 216
rect 487 199 504 216
rect 521 199 538 216
rect 555 199 572 216
rect 589 199 606 216
rect 623 199 640 216
rect 657 199 674 216
rect 691 199 708 216
rect 725 199 742 216
rect 759 199 776 216
rect 793 199 810 216
rect 827 199 844 216
rect 861 199 878 216
rect 895 199 912 216
rect 929 199 946 216
rect 963 204 1067 216
rect 1084 204 1096 221
rect 963 199 1096 204
rect 462 198 1096 199
rect 265 166 431 174
rect 265 146 408 166
rect 429 146 431 166
rect 462 168 1115 169
rect 462 151 470 168
rect 487 151 504 168
rect 521 151 538 168
rect 555 151 572 168
rect 589 151 606 168
rect 623 151 640 168
rect 657 151 674 168
rect 691 151 708 168
rect 725 151 742 168
rect 759 151 776 168
rect 793 151 810 168
rect 827 151 844 168
rect 861 151 878 168
rect 895 151 912 168
rect 929 151 946 168
rect 963 151 1115 168
rect 462 150 1115 151
rect 141 124 142 141
rect 159 124 160 141
rect 141 107 160 124
rect 141 90 142 107
rect 159 90 160 107
rect 141 73 160 90
rect 217 129 236 146
rect 217 112 218 129
rect 235 112 236 129
rect 217 95 236 112
rect 217 78 218 95
rect 235 78 236 95
rect 217 70 236 78
rect 265 142 431 146
rect 265 125 266 142
rect 283 138 431 142
rect 283 125 284 138
rect 265 108 284 125
rect 1017 110 1042 150
rect 1060 146 1115 150
rect 1067 142 1115 146
rect 1072 137 1115 142
rect 1073 134 1115 137
rect 1073 117 1086 134
rect 1103 117 1115 134
rect 265 91 266 108
rect 283 91 284 108
rect 1013 93 1021 110
rect 1038 93 1046 110
rect 265 74 284 91
rect 1073 89 1115 90
rect 322 67 390 73
rect 1073 69 1086 89
rect 1103 69 1115 89
rect 1160 78 1241 82
rect 322 50 343 67
rect 360 50 390 67
rect 322 32 390 50
rect 1160 61 1180 78
rect 1197 61 1241 78
rect 1160 32 1241 61
rect 0 15 21 32
rect 38 15 55 32
rect 72 15 89 32
rect 106 15 123 32
rect 140 15 157 32
rect 174 15 191 32
rect 208 15 225 32
rect 242 15 259 32
rect 276 15 293 32
rect 310 15 327 32
rect 344 15 361 32
rect 378 15 395 32
rect 412 15 429 32
rect 446 15 463 32
rect 480 15 497 32
rect 514 15 531 32
rect 548 15 565 32
rect 582 15 599 32
rect 616 15 633 32
rect 650 15 667 32
rect 684 15 701 32
rect 718 15 735 32
rect 752 15 769 32
rect 786 15 803 32
rect 820 15 837 32
rect 854 15 871 32
rect 888 15 905 32
rect 922 15 939 32
rect 956 15 973 32
rect 990 15 1007 32
rect 1024 15 1041 32
rect 1058 15 1075 32
rect 1092 15 1109 32
rect 1126 15 1143 32
rect 1160 15 1177 32
rect 1194 15 1211 32
rect 1228 15 1245 32
rect 1262 15 1279 32
rect 1296 15 1313 32
rect 1330 15 1347 32
rect 1364 15 1381 32
rect 1398 15 1415 32
rect 1432 15 1449 32
rect 1466 15 1483 32
rect 1500 15 1517 32
rect 1534 15 1551 32
rect 1568 15 1585 32
rect 1602 15 1619 32
rect 1636 15 1653 32
rect 1670 15 1687 32
rect 1704 15 1721 32
rect 1738 15 1755 32
rect 1772 15 1789 32
rect 1806 15 1823 32
rect 1840 15 1857 32
rect 1874 15 1891 32
rect 1908 15 1925 32
rect 1942 15 1959 32
rect 1976 15 1993 32
rect 2010 15 2067 32
<< viali >>
rect 21 607 38 624
rect 55 607 72 624
rect 89 607 106 624
rect 123 607 140 624
rect 157 607 174 624
rect 191 607 208 624
rect 225 607 242 624
rect 259 607 276 624
rect 293 607 310 624
rect 327 607 344 624
rect 361 607 378 624
rect 395 607 412 624
rect 429 607 446 624
rect 463 607 480 624
rect 497 607 514 624
rect 531 607 548 624
rect 565 607 582 624
rect 599 607 616 624
rect 633 607 650 624
rect 667 607 684 624
rect 701 607 718 624
rect 735 607 752 624
rect 769 607 786 624
rect 803 607 820 624
rect 837 607 854 624
rect 871 607 888 624
rect 905 607 922 624
rect 939 607 956 624
rect 973 607 990 624
rect 1007 607 1024 624
rect 1041 607 1058 624
rect 1075 607 1092 624
rect 1109 607 1126 624
rect 1143 607 1160 624
rect 1177 607 1194 624
rect 1211 607 1228 624
rect 1245 607 1262 624
rect 1279 607 1296 624
rect 1313 607 1330 624
rect 1347 607 1364 624
rect 1381 607 1398 624
rect 1415 607 1432 624
rect 1449 607 1466 624
rect 1483 607 1500 624
rect 1517 607 1534 624
rect 1551 607 1568 624
rect 1585 607 1602 624
rect 1619 607 1636 624
rect 1653 607 1670 624
rect 1687 607 1704 624
rect 1721 607 1738 624
rect 1755 607 1772 624
rect 1789 607 1806 624
rect 1823 607 1840 624
rect 1857 607 1874 624
rect 1891 607 1908 624
rect 1925 607 1942 624
rect 1959 607 1976 624
rect 1993 607 2010 624
rect 2027 607 2044 624
rect 1281 540 1294 557
rect 1294 540 1298 557
rect 1315 540 1328 557
rect 1328 540 1332 557
rect 204 411 221 428
rect 1130 408 1147 425
rect 1882 422 1899 439
rect 1925 422 1942 439
rect 21 310 38 327
rect 55 310 72 327
rect 89 310 106 327
rect 123 310 140 327
rect 157 310 174 327
rect 191 310 208 327
rect 225 310 242 327
rect 259 310 276 327
rect 293 310 310 327
rect 327 310 344 327
rect 361 310 378 327
rect 395 310 412 327
rect 429 310 446 327
rect 463 310 480 327
rect 497 310 514 327
rect 531 310 548 327
rect 565 310 582 327
rect 599 310 616 327
rect 633 310 650 327
rect 667 310 684 327
rect 701 310 718 327
rect 735 310 752 327
rect 769 310 786 327
rect 803 310 820 327
rect 837 310 854 327
rect 871 310 888 327
rect 905 310 922 327
rect 939 310 956 327
rect 973 310 990 327
rect 1007 310 1024 327
rect 146 254 163 271
rect 78 166 95 183
rect 94 111 111 128
rect 94 77 111 94
rect 1010 257 1027 274
rect 1143 310 1160 327
rect 1177 310 1194 327
rect 1211 310 1228 327
rect 1245 310 1262 327
rect 1279 310 1296 327
rect 1313 310 1330 327
rect 1347 310 1364 327
rect 1381 310 1398 327
rect 1415 310 1432 327
rect 1449 310 1466 327
rect 1483 310 1500 327
rect 1517 310 1534 327
rect 1551 310 1568 327
rect 1585 310 1602 327
rect 1619 310 1636 327
rect 1653 310 1670 327
rect 1687 310 1704 327
rect 1721 310 1738 327
rect 1755 310 1772 327
rect 1789 310 1806 327
rect 1823 310 1840 327
rect 1857 310 1874 327
rect 1891 310 1908 327
rect 1925 310 1942 327
rect 1959 310 1976 327
rect 1993 310 2010 327
rect 202 166 219 183
rect 218 112 235 129
rect 218 78 235 95
rect 1086 86 1103 89
rect 1086 72 1103 86
rect 21 15 38 32
rect 55 15 72 32
rect 89 15 106 32
rect 123 15 140 32
rect 157 15 174 32
rect 191 15 208 32
rect 225 15 242 32
rect 259 15 276 32
rect 293 15 310 32
rect 327 15 344 32
rect 361 15 378 32
rect 395 15 412 32
rect 429 15 446 32
rect 463 15 480 32
rect 497 15 514 32
rect 531 15 548 32
rect 565 15 582 32
rect 599 15 616 32
rect 633 15 650 32
rect 667 15 684 32
rect 701 15 718 32
rect 735 15 752 32
rect 769 15 786 32
rect 803 15 820 32
rect 837 15 854 32
rect 871 15 888 32
rect 905 15 922 32
rect 939 15 956 32
rect 973 15 990 32
rect 1007 15 1024 32
rect 1041 15 1058 32
rect 1075 15 1092 32
rect 1109 15 1126 32
rect 1143 15 1160 32
rect 1177 15 1194 32
rect 1211 15 1228 32
rect 1245 15 1262 32
rect 1279 15 1296 32
rect 1313 15 1330 32
rect 1347 15 1364 32
rect 1381 15 1398 32
rect 1415 15 1432 32
rect 1449 15 1466 32
rect 1483 15 1500 32
rect 1517 15 1534 32
rect 1551 15 1568 32
rect 1585 15 1602 32
rect 1619 15 1636 32
rect 1653 15 1670 32
rect 1687 15 1704 32
rect 1721 15 1738 32
rect 1755 15 1772 32
rect 1789 15 1806 32
rect 1823 15 1840 32
rect 1857 15 1874 32
rect 1891 15 1908 32
rect 1925 15 1942 32
rect 1959 15 1976 32
rect 1993 15 2010 32
<< metal1 >>
rect 0 624 2066 640
rect 0 607 21 624
rect 38 607 55 624
rect 72 607 89 624
rect 106 607 123 624
rect 140 607 157 624
rect 174 607 191 624
rect 208 607 225 624
rect 242 607 259 624
rect 276 607 293 624
rect 310 607 327 624
rect 344 607 361 624
rect 378 607 395 624
rect 412 607 429 624
rect 446 607 463 624
rect 480 607 497 624
rect 514 607 531 624
rect 548 607 565 624
rect 582 607 599 624
rect 616 607 633 624
rect 650 607 667 624
rect 684 607 701 624
rect 718 607 735 624
rect 752 607 769 624
rect 786 607 803 624
rect 820 607 837 624
rect 854 607 871 624
rect 888 607 905 624
rect 922 607 939 624
rect 956 607 973 624
rect 990 607 1007 624
rect 1024 607 1041 624
rect 1058 607 1075 624
rect 1092 607 1109 624
rect 1126 607 1143 624
rect 1160 607 1177 624
rect 1194 607 1211 624
rect 1228 607 1245 624
rect 1262 607 1279 624
rect 1296 607 1313 624
rect 1330 607 1347 624
rect 1364 607 1381 624
rect 1398 607 1415 624
rect 1432 607 1449 624
rect 1466 607 1483 624
rect 1500 607 1517 624
rect 1534 607 1551 624
rect 1568 607 1585 624
rect 1602 607 1619 624
rect 1636 607 1653 624
rect 1670 607 1687 624
rect 1704 607 1721 624
rect 1738 607 1755 624
rect 1772 607 1789 624
rect 1806 607 1823 624
rect 1840 607 1857 624
rect 1874 607 1891 624
rect 1908 607 1925 624
rect 1942 607 1959 624
rect 1976 607 1993 624
rect 2010 607 2027 624
rect 2044 607 2066 624
rect 0 592 2066 607
rect 1275 560 1343 563
rect 1275 557 1293 560
rect 1319 557 1343 560
rect 1275 540 1281 557
rect 1332 540 1343 557
rect 1275 534 1293 540
rect 1319 534 1343 540
rect 1876 446 1946 592
rect 1876 439 1948 446
rect 196 432 228 435
rect 196 406 199 432
rect 225 406 228 432
rect 196 403 228 406
rect 1122 429 1154 432
rect 1122 403 1125 429
rect 1151 403 1154 429
rect 1876 422 1882 439
rect 1899 422 1925 439
rect 1942 422 1948 439
rect 1876 416 1948 422
rect 1122 402 1154 403
rect 1 327 2066 344
rect 1 310 21 327
rect 38 310 55 327
rect 72 310 89 327
rect 106 310 123 327
rect 140 310 157 327
rect 174 310 191 327
rect 208 310 225 327
rect 242 310 259 327
rect 276 310 293 327
rect 310 310 327 327
rect 344 310 361 327
rect 378 310 395 327
rect 412 310 429 327
rect 446 310 463 327
rect 480 310 497 327
rect 514 310 531 327
rect 548 310 565 327
rect 582 310 599 327
rect 616 310 633 327
rect 650 310 667 327
rect 684 310 701 327
rect 718 310 735 327
rect 752 310 769 327
rect 786 310 803 327
rect 820 310 837 327
rect 854 310 871 327
rect 888 310 905 327
rect 922 310 939 327
rect 956 310 973 327
rect 990 310 1007 327
rect 1024 310 1143 327
rect 1160 310 1177 327
rect 1194 310 1211 327
rect 1228 310 1245 327
rect 1262 310 1279 327
rect 1296 310 1313 327
rect 1330 310 1347 327
rect 1364 310 1381 327
rect 1398 310 1415 327
rect 1432 310 1449 327
rect 1466 310 1483 327
rect 1500 310 1517 327
rect 1534 310 1551 327
rect 1568 310 1585 327
rect 1602 310 1619 327
rect 1636 310 1653 327
rect 1670 310 1687 327
rect 1704 310 1721 327
rect 1738 310 1755 327
rect 1772 310 1789 327
rect 1806 310 1823 327
rect 1840 310 1857 327
rect 1874 310 1891 327
rect 1908 310 1925 327
rect 1942 310 1959 327
rect 1976 310 1993 327
rect 2010 310 2066 327
rect 1 296 2066 310
rect 1002 278 1034 281
rect 138 275 170 278
rect 138 249 141 275
rect 167 249 170 275
rect 1002 252 1005 278
rect 1031 252 1034 278
rect 1002 249 1034 252
rect 138 246 170 249
rect 1268 210 1347 229
rect 71 187 103 190
rect 71 161 74 187
rect 100 161 103 187
rect 71 158 103 161
rect 194 187 226 190
rect 194 161 197 187
rect 223 161 226 187
rect 194 158 226 161
rect 1268 174 1281 210
rect 1335 174 1347 210
rect 1268 154 1347 174
rect 90 128 115 134
rect 90 111 94 128
rect 111 111 115 128
rect 90 99 115 111
rect 214 129 239 135
rect 214 112 218 129
rect 235 112 239 129
rect 214 99 239 112
rect 1268 99 1316 154
rect 90 95 1316 99
rect 90 94 218 95
rect 90 77 94 94
rect 111 78 218 94
rect 235 89 1316 95
rect 235 78 1086 89
rect 111 77 1086 78
rect 90 72 1086 77
rect 1103 72 1316 89
rect 90 69 1316 72
rect 0 32 2067 48
rect 0 15 21 32
rect 38 15 55 32
rect 72 15 89 32
rect 106 15 123 32
rect 140 15 157 32
rect 174 15 191 32
rect 208 15 225 32
rect 242 15 259 32
rect 276 15 293 32
rect 310 15 327 32
rect 344 15 361 32
rect 378 15 395 32
rect 412 15 429 32
rect 446 15 463 32
rect 480 15 497 32
rect 514 15 531 32
rect 548 15 565 32
rect 582 15 599 32
rect 616 15 633 32
rect 650 15 667 32
rect 684 15 701 32
rect 718 15 735 32
rect 752 15 769 32
rect 786 15 803 32
rect 820 15 837 32
rect 854 15 871 32
rect 888 15 905 32
rect 922 15 939 32
rect 956 15 973 32
rect 990 15 1007 32
rect 1024 15 1041 32
rect 1058 15 1075 32
rect 1092 15 1109 32
rect 1126 15 1143 32
rect 1160 15 1177 32
rect 1194 15 1211 32
rect 1228 15 1245 32
rect 1262 15 1279 32
rect 1296 15 1313 32
rect 1330 15 1347 32
rect 1364 15 1381 32
rect 1398 15 1415 32
rect 1432 15 1449 32
rect 1466 15 1483 32
rect 1500 15 1517 32
rect 1534 15 1551 32
rect 1568 15 1585 32
rect 1602 15 1619 32
rect 1636 15 1653 32
rect 1670 15 1687 32
rect 1704 15 1721 32
rect 1738 15 1755 32
rect 1772 15 1789 32
rect 1806 15 1823 32
rect 1840 15 1857 32
rect 1874 15 1891 32
rect 1908 15 1925 32
rect 1942 15 1959 32
rect 1976 15 1993 32
rect 2010 15 2067 32
rect 0 0 2067 15
<< via1 >>
rect 1293 557 1319 560
rect 1293 540 1298 557
rect 1298 540 1315 557
rect 1315 540 1319 557
rect 1293 534 1319 540
rect 199 428 225 432
rect 199 411 204 428
rect 204 411 221 428
rect 221 411 225 428
rect 199 406 225 411
rect 1125 425 1151 429
rect 1125 408 1130 425
rect 1130 408 1147 425
rect 1147 408 1151 425
rect 1125 403 1151 408
rect 141 271 167 275
rect 141 254 146 271
rect 146 254 163 271
rect 163 254 167 271
rect 141 249 167 254
rect 1005 274 1031 278
rect 1005 257 1010 274
rect 1010 257 1027 274
rect 1027 257 1031 274
rect 1005 252 1031 257
rect 74 183 100 187
rect 74 166 78 183
rect 78 166 95 183
rect 95 166 100 183
rect 74 161 100 166
rect 197 183 223 187
rect 197 166 202 183
rect 202 166 219 183
rect 219 166 223 183
rect 197 161 223 166
rect 1281 174 1335 210
<< metal2 >>
rect 1278 560 1339 563
rect 1278 534 1293 560
rect 1319 534 1339 560
rect 184 433 228 435
rect 60 432 228 433
rect 60 406 199 432
rect 225 406 228 432
rect 60 403 228 406
rect 870 429 1154 432
rect 870 403 1125 429
rect 1151 403 1154 429
rect 60 397 227 403
rect 870 400 1154 403
rect 60 272 92 397
rect 870 300 917 400
rect 1 241 92 272
rect 138 275 917 300
rect 138 249 141 275
rect 167 260 917 275
rect 947 278 1034 281
rect 167 249 170 260
rect 138 246 170 249
rect 947 252 1005 278
rect 1031 252 1034 278
rect 947 249 1034 252
rect 60 190 92 241
rect 60 187 103 190
rect 60 161 74 187
rect 100 161 103 187
rect 60 158 103 161
rect 176 187 226 190
rect 176 161 197 187
rect 223 161 226 187
rect 176 110 209 161
rect 947 110 984 249
rect 1278 210 1339 534
rect 1278 174 1281 210
rect 1335 174 1339 210
rect 1278 171 1339 174
rect 176 109 984 110
rect 1 73 984 109
<< labels >>
rlabel metal1 0 592 0 640 3 VDD
port 1 e power bidirectional
rlabel metal1 1 296 1 344 3 GND
port 2 e ground bidirectional
rlabel metal1 0 0 0 48 3 VDD
port 1 e power bidirectional
rlabel metal2 1 73 1 109 3 Up
port 3 e signal input
rlabel metal2 1 241 1 272 3 Down
port 4 e signal input
rlabel locali 2066 349 2066 402 7 Out
port 5 w signal output
rlabel locali 51 481 51 505 3 ENb
port 6 e signal input
<< properties >>
string LEFclass CORE
string LEFsite unithddb1
<< end >>
