magic
tech sky130A
timestamp 1605926473
<< nwell >>
rect 0 185 932 320
rect 0 149 237 185
rect 396 184 932 185
rect 396 149 510 184
rect 667 160 932 184
rect 667 155 786 160
rect 679 148 786 155
<< nmos >>
rect 64 75 79 111
rect 175 75 190 111
rect 317 67 332 151
rect 448 74 463 110
rect 582 66 597 150
rect 714 75 729 111
rect 818 62 833 98
rect 869 62 884 98
<< pmos >>
rect 64 173 79 245
rect 175 173 190 245
rect 317 204 332 246
rect 448 172 463 244
rect 582 203 597 245
rect 714 173 729 245
rect 818 183 833 255
rect 869 183 884 255
<< ndiff >>
rect 288 142 317 151
rect 288 125 294 142
rect 311 125 317 142
rect 35 102 64 111
rect 35 85 41 102
rect 58 85 64 102
rect 35 75 64 85
rect 79 102 108 111
rect 79 85 85 102
rect 102 85 108 102
rect 79 75 108 85
rect 146 102 175 111
rect 146 85 152 102
rect 169 85 175 102
rect 146 75 175 85
rect 190 102 219 111
rect 190 85 196 102
rect 213 85 219 102
rect 288 108 317 125
rect 190 75 219 85
rect 288 91 294 108
rect 311 91 317 108
rect 288 67 317 91
rect 332 142 361 151
rect 332 125 338 142
rect 355 125 361 142
rect 332 108 361 125
rect 553 141 582 150
rect 553 124 559 141
rect 576 124 582 141
rect 332 91 338 108
rect 355 91 361 108
rect 332 67 361 91
rect 419 101 448 110
rect 419 84 425 101
rect 442 84 448 101
rect 419 74 448 84
rect 463 101 492 110
rect 463 84 469 101
rect 486 84 492 101
rect 553 107 582 124
rect 463 74 492 84
rect 553 90 559 107
rect 576 90 582 107
rect 553 66 582 90
rect 597 141 626 150
rect 597 124 603 141
rect 620 124 626 141
rect 597 107 626 124
rect 597 90 603 107
rect 620 90 626 107
rect 597 66 626 90
rect 685 102 714 111
rect 685 85 691 102
rect 708 85 714 102
rect 685 75 714 85
rect 729 102 758 111
rect 729 85 735 102
rect 752 85 758 102
rect 729 75 758 85
rect 787 88 818 98
rect 787 71 793 88
rect 810 71 818 88
rect 787 62 818 71
rect 833 83 869 98
rect 833 66 845 83
rect 862 66 869 83
rect 833 62 869 66
rect 884 88 913 98
rect 884 71 892 88
rect 909 71 913 88
rect 884 62 913 71
<< pdiff >>
rect 35 241 64 245
rect 35 224 41 241
rect 58 224 64 241
rect 35 207 64 224
rect 35 190 41 207
rect 58 190 64 207
rect 35 173 64 190
rect 79 228 108 245
rect 79 211 85 228
rect 102 211 108 228
rect 79 194 108 211
rect 79 177 85 194
rect 102 177 108 194
rect 79 173 108 177
rect 146 241 175 245
rect 146 224 152 241
rect 169 224 175 241
rect 146 207 175 224
rect 146 190 152 207
rect 169 190 175 207
rect 146 173 175 190
rect 190 228 219 245
rect 190 211 196 228
rect 213 211 219 228
rect 288 233 317 246
rect 190 194 219 211
rect 288 216 294 233
rect 311 216 317 233
rect 288 204 317 216
rect 332 232 361 246
rect 332 215 338 232
rect 355 215 361 232
rect 332 204 361 215
rect 419 240 448 244
rect 419 223 425 240
rect 442 223 448 240
rect 419 206 448 223
rect 190 177 196 194
rect 213 177 219 194
rect 190 173 219 177
rect 419 189 425 206
rect 442 189 448 206
rect 419 172 448 189
rect 463 227 492 244
rect 463 210 469 227
rect 486 210 492 227
rect 463 193 492 210
rect 553 232 582 245
rect 553 215 559 232
rect 576 215 582 232
rect 553 203 582 215
rect 597 231 626 245
rect 597 214 603 231
rect 620 214 626 231
rect 787 251 818 255
rect 685 241 714 245
rect 685 224 691 241
rect 708 224 714 241
rect 597 203 626 214
rect 685 207 714 224
rect 463 176 469 193
rect 486 176 492 193
rect 685 190 691 207
rect 708 190 714 207
rect 463 172 492 176
rect 685 173 714 190
rect 729 228 758 245
rect 729 211 735 228
rect 752 211 758 228
rect 729 194 758 211
rect 729 177 735 194
rect 752 177 758 194
rect 787 234 793 251
rect 810 234 818 251
rect 787 217 818 234
rect 787 200 793 217
rect 810 200 818 217
rect 787 183 818 200
rect 833 251 869 255
rect 833 234 844 251
rect 861 234 869 251
rect 833 183 869 234
rect 884 251 914 255
rect 884 234 891 251
rect 908 234 914 251
rect 884 217 914 234
rect 884 200 891 217
rect 908 200 914 217
rect 884 183 913 200
rect 729 173 758 177
<< ndiffc >>
rect 294 125 311 142
rect 41 85 58 102
rect 85 85 102 102
rect 152 85 169 102
rect 196 85 213 102
rect 294 91 311 108
rect 338 125 355 142
rect 559 124 576 141
rect 338 91 355 108
rect 425 84 442 101
rect 469 84 486 101
rect 559 90 576 107
rect 603 124 620 141
rect 603 90 620 107
rect 691 85 708 102
rect 735 85 752 102
rect 793 71 810 88
rect 845 66 862 83
rect 892 71 909 88
<< pdiffc >>
rect 41 224 58 241
rect 41 190 58 207
rect 85 211 102 228
rect 85 177 102 194
rect 152 224 169 241
rect 152 190 169 207
rect 196 211 213 228
rect 294 216 311 233
rect 338 215 355 232
rect 425 223 442 240
rect 196 177 213 194
rect 425 189 442 206
rect 469 210 486 227
rect 559 215 576 232
rect 603 214 620 231
rect 691 224 708 241
rect 469 176 486 193
rect 691 190 708 207
rect 735 211 752 228
rect 735 177 752 194
rect 793 234 810 251
rect 793 200 810 217
rect 844 234 861 251
rect 891 234 908 251
rect 891 200 908 217
<< psubdiff >>
rect 3 15 16 32
rect 33 15 45 32
rect 87 15 100 32
rect 117 15 129 32
rect 167 15 180 32
rect 197 15 209 32
rect 302 15 315 32
rect 332 15 344 32
rect 394 15 407 32
rect 424 15 436 32
rect 500 15 513 32
rect 530 15 542 32
rect 584 15 597 32
rect 614 15 626 32
rect 702 15 715 32
rect 732 15 744 32
rect 786 15 799 32
rect 816 15 828 32
rect 870 15 883 32
rect 900 15 912 32
<< nsubdiff >>
rect 43 283 55 302
rect 74 283 86 302
rect 125 283 137 302
rect 156 283 168 302
rect 270 283 282 302
rect 301 283 313 302
rect 348 283 360 302
rect 379 283 391 302
rect 442 283 454 302
rect 473 283 485 302
rect 550 283 562 302
rect 581 283 593 302
rect 670 283 682 302
rect 701 283 713 302
rect 756 283 768 302
rect 787 283 799 302
rect 842 283 854 302
rect 873 283 885 302
<< psubdiffcont >>
rect 16 15 33 32
rect 100 15 117 32
rect 180 15 197 32
rect 315 15 332 32
rect 407 15 424 32
rect 513 15 530 32
rect 597 15 614 32
rect 715 15 732 32
rect 799 15 816 32
rect 883 15 900 32
<< nsubdiffcont >>
rect 55 283 74 302
rect 137 283 156 302
rect 282 283 301 302
rect 360 283 379 302
rect 454 283 473 302
rect 562 283 581 302
rect 682 283 701 302
rect 768 283 787 302
rect 854 283 873 302
<< poly >>
rect 64 245 79 258
rect 175 245 190 258
rect 239 257 332 272
rect 239 247 266 257
rect 239 230 244 247
rect 261 230 266 247
rect 317 246 332 257
rect 239 222 266 230
rect 448 244 463 257
rect 582 256 671 271
rect 582 245 597 256
rect 317 190 332 204
rect 64 153 79 173
rect 175 153 190 173
rect 644 241 671 256
rect 714 245 729 258
rect 818 255 833 268
rect 869 255 884 268
rect 644 224 649 241
rect 666 224 671 241
rect 644 216 671 224
rect 582 189 597 203
rect 35 151 79 153
rect 146 151 190 153
rect 317 151 332 164
rect 448 152 463 172
rect 32 148 79 151
rect 32 131 41 148
rect 58 131 79 148
rect 32 127 79 131
rect 143 148 190 151
rect 143 131 152 148
rect 169 131 190 148
rect 143 127 190 131
rect 35 126 79 127
rect 146 126 190 127
rect 64 111 79 126
rect 175 111 190 126
rect 240 92 267 100
rect 240 75 245 92
rect 262 75 267 92
rect 64 62 79 75
rect 175 62 190 75
rect 240 59 267 75
rect 419 150 463 152
rect 582 150 597 163
rect 714 153 729 173
rect 818 164 833 183
rect 869 168 884 183
rect 866 164 884 168
rect 805 159 833 164
rect 685 151 729 153
rect 416 147 463 150
rect 416 130 425 147
rect 442 130 463 147
rect 416 126 463 130
rect 419 125 463 126
rect 448 110 463 125
rect 512 88 539 96
rect 317 59 332 67
rect 448 61 463 74
rect 512 71 517 88
rect 534 71 539 88
rect 240 44 332 59
rect 512 58 539 71
rect 682 148 729 151
rect 682 131 691 148
rect 708 131 729 148
rect 802 142 810 159
rect 827 142 834 159
rect 855 155 884 164
rect 805 137 833 142
rect 682 127 729 131
rect 685 126 729 127
rect 714 111 729 126
rect 818 98 833 137
rect 855 138 860 155
rect 877 138 884 155
rect 855 130 884 138
rect 866 124 884 130
rect 869 98 884 124
rect 582 58 597 66
rect 714 62 729 75
rect 512 43 597 58
rect 818 49 833 62
rect 869 49 884 62
<< polycont >>
rect 244 230 261 247
rect 649 224 666 241
rect 41 131 58 148
rect 152 131 169 148
rect 245 75 262 92
rect 425 130 442 147
rect 517 71 534 88
rect 691 131 708 148
rect 810 142 827 159
rect 860 138 877 155
<< locali >>
rect 0 283 55 302
rect 74 283 137 302
rect 156 283 282 302
rect 301 283 360 302
rect 379 283 454 302
rect 473 283 562 302
rect 581 283 682 302
rect 701 283 768 302
rect 787 283 854 302
rect 873 283 932 302
rect 41 241 58 283
rect 41 207 58 224
rect 41 173 58 190
rect 85 228 102 245
rect 85 194 102 211
rect 85 156 102 177
rect 152 241 169 283
rect 244 247 261 255
rect 152 207 169 224
rect 152 173 169 190
rect 196 228 213 245
rect 244 222 261 229
rect 294 233 311 246
rect 196 194 213 211
rect 294 193 311 216
rect 196 157 213 177
rect 239 163 311 193
rect 239 157 264 163
rect 85 149 115 156
rect 0 131 41 148
rect 58 131 66 148
rect 85 132 91 149
rect 108 132 115 149
rect 85 126 115 132
rect 143 131 152 148
rect 169 131 177 148
rect 196 127 264 157
rect 294 142 311 163
rect 41 102 58 111
rect 41 32 58 85
rect 85 102 102 126
rect 85 75 102 85
rect 152 102 169 111
rect 152 32 169 85
rect 196 102 213 127
rect 294 108 311 125
rect 196 75 213 85
rect 237 75 245 92
rect 262 75 270 92
rect 294 83 311 91
rect 338 232 355 246
rect 338 190 355 215
rect 425 240 442 283
rect 425 206 442 223
rect 338 163 408 190
rect 425 172 442 189
rect 469 227 486 244
rect 469 193 486 210
rect 559 232 576 245
rect 559 191 576 215
rect 338 142 355 163
rect 391 154 408 163
rect 469 156 486 176
rect 509 162 576 191
rect 509 156 537 162
rect 391 152 412 154
rect 391 147 446 152
rect 391 130 425 147
rect 442 130 450 147
rect 391 127 446 130
rect 469 127 537 156
rect 559 141 576 162
rect 338 108 355 125
rect 338 83 355 91
rect 425 101 442 110
rect 237 74 270 75
rect 425 32 442 84
rect 469 101 486 127
rect 559 107 576 124
rect 469 74 486 84
rect 509 71 517 88
rect 534 71 542 88
rect 559 82 576 90
rect 603 231 620 245
rect 649 241 666 250
rect 649 216 666 224
rect 691 241 708 283
rect 790 251 812 259
rect 603 188 620 214
rect 691 207 708 224
rect 603 163 657 188
rect 691 173 708 190
rect 735 228 752 245
rect 735 194 752 211
rect 790 234 793 251
rect 810 234 812 251
rect 790 217 812 234
rect 841 251 864 283
rect 841 234 844 251
rect 861 234 864 251
rect 841 222 864 234
rect 891 255 909 259
rect 891 251 920 255
rect 908 234 920 251
rect 790 200 793 217
rect 810 201 812 217
rect 891 217 920 234
rect 810 200 874 201
rect 790 184 874 200
rect 603 141 620 163
rect 603 107 620 124
rect 603 82 620 90
rect 638 152 657 163
rect 735 156 752 177
rect 855 164 874 184
rect 908 200 920 217
rect 891 181 920 200
rect 895 164 920 181
rect 679 152 712 153
rect 638 148 712 152
rect 735 149 769 156
rect 638 131 691 148
rect 708 131 716 148
rect 735 132 744 149
rect 761 132 769 149
rect 801 142 810 159
rect 827 142 835 159
rect 855 155 877 164
rect 855 138 860 155
rect 855 135 877 138
rect 638 128 712 131
rect 638 101 657 128
rect 735 126 769 132
rect 854 130 877 135
rect 691 102 708 111
rect 638 94 666 101
rect 638 77 646 94
rect 663 77 666 94
rect 638 70 666 77
rect 691 32 708 85
rect 735 102 752 126
rect 854 125 872 130
rect 735 75 752 85
rect 789 108 872 125
rect 789 88 811 108
rect 903 98 920 164
rect 789 71 793 88
rect 810 71 811 88
rect 789 62 811 71
rect 842 83 864 91
rect 842 66 845 83
rect 862 66 864 83
rect 842 32 864 66
rect 890 88 920 98
rect 890 71 892 88
rect 909 71 920 88
rect 890 62 920 71
rect 0 15 16 32
rect 33 15 100 32
rect 117 15 180 32
rect 197 15 315 32
rect 332 15 407 32
rect 424 15 513 32
rect 530 15 597 32
rect 614 15 715 32
rect 732 15 799 32
rect 816 15 883 32
rect 900 15 935 32
<< viali >>
rect 55 283 74 302
rect 137 283 156 302
rect 282 283 301 302
rect 360 283 379 302
rect 454 283 473 302
rect 562 283 581 302
rect 682 283 701 302
rect 768 283 787 302
rect 854 283 873 302
rect 244 230 261 247
rect 244 229 261 230
rect 41 131 58 148
rect 91 132 108 149
rect 152 131 169 148
rect 245 75 262 92
rect 517 71 534 88
rect 649 224 666 241
rect 744 132 761 149
rect 810 142 827 159
rect 646 77 663 94
rect 16 15 33 32
rect 100 15 117 32
rect 180 15 197 32
rect 315 15 332 32
rect 407 15 424 32
rect 513 15 530 32
rect 597 15 614 32
rect 715 15 732 32
rect 799 15 816 32
rect 883 15 900 32
<< metal1 >>
rect 0 302 932 320
rect 0 283 55 302
rect 74 283 137 302
rect 156 283 282 302
rect 301 283 360 302
rect 379 283 454 302
rect 473 283 562 302
rect 581 283 682 302
rect 701 283 768 302
rect 787 283 854 302
rect 873 283 932 302
rect 0 272 932 283
rect 237 251 269 254
rect 35 218 157 250
rect 237 225 240 251
rect 266 225 269 251
rect 644 249 672 250
rect 237 222 269 225
rect 643 241 672 249
rect 643 224 649 241
rect 666 224 672 241
rect 35 148 64 218
rect 132 207 157 218
rect 643 207 672 224
rect 132 182 672 207
rect 804 159 835 165
rect 35 131 41 148
rect 58 131 64 148
rect 35 127 64 131
rect 36 98 64 127
rect 83 155 118 159
rect 83 129 88 155
rect 114 129 118 155
rect 83 124 118 129
rect 146 149 769 154
rect 146 148 744 149
rect 146 131 152 148
rect 169 132 744 148
rect 761 132 769 149
rect 804 142 810 159
rect 827 142 835 159
rect 804 137 835 142
rect 169 131 769 132
rect 146 126 769 131
rect 807 100 834 137
rect 36 92 271 98
rect 36 75 245 92
rect 262 75 271 92
rect 36 69 271 75
rect 508 93 541 96
rect 508 66 511 93
rect 538 66 541 93
rect 640 94 834 100
rect 640 77 646 94
rect 663 77 834 94
rect 640 73 834 77
rect 640 71 672 73
rect 641 70 672 71
rect 508 63 541 66
rect 0 32 935 48
rect 0 15 16 32
rect 33 15 100 32
rect 117 15 180 32
rect 197 15 315 32
rect 332 15 407 32
rect 424 15 513 32
rect 530 15 597 32
rect 614 15 715 32
rect 732 15 799 32
rect 816 15 883 32
rect 900 15 935 32
rect 0 0 935 15
<< via1 >>
rect 240 247 266 251
rect 240 229 244 247
rect 244 229 261 247
rect 261 229 266 247
rect 240 225 266 229
rect 88 149 114 155
rect 88 132 91 149
rect 91 132 108 149
rect 108 132 114 149
rect 88 129 114 132
rect 511 88 538 93
rect 511 71 517 88
rect 517 71 534 88
rect 534 71 538 88
rect 511 66 538 71
<< metal2 >>
rect 237 225 240 251
rect 266 225 269 251
rect 85 159 118 166
rect 83 157 118 159
rect 237 157 269 225
rect 83 155 540 157
rect 83 129 88 155
rect 114 129 540 155
rect 83 128 540 129
rect 83 124 118 128
rect 507 93 540 128
rect 507 87 511 93
rect 508 66 511 87
rect 538 66 541 93
rect 508 63 541 66
<< labels >>
rlabel locali 905 138 919 152 1 Clk_Out
port 3 n
rlabel locali 0 131 0 148 3 Clk_In
port 5 e
rlabel metal1 0 0 0 48 3 GND
port 4 e
rlabel metal1 0 272 0 320 3 VDD
port 6 e
<< properties >>
string LEFsite unithddb1
string LEFclass CORE
<< end >>
